PK   -�eTv��#  h�     cirkitFile.json�]���6����g")~����pm��h�%QY�{O����<н�=ӑ�wmˢ5�p�A�E�G���O���G��h�bY��G[�f��膰�����'sx6��g��z9}_�����g����I��p�\��z�*#�L��
�%Y�Mb�	I%�"+�,�4ݼ�XY�W��	c�$Yii�e.�B��q͋�Hw�������n�AS��)Fj���=�Z3��Bj��:�H�R3��#�@H�a��%Bj��Zb�V�Fj�kͩ����9I��ʪ�p�&e%5+�yjݵ�5����(m$�9b��)�S���]hl��<M���*�4�Z�2W�jH��@����� mJ9H��Rʪ�Ieswע���V'�ɩ������rS�Z&�LU��H�I*+[�*���5n��-�����,J757*ɕ�i�-Tɫ���!#�֚����ݹ�ZX�-�D��T�TZh�{"!jfT𩻍Yn�,rÒT	�^���%O4���y!��E����$h`�3u(���]�t1J������-BjL��1R��*� ]�q�D�%�SD�(��x̂�$��!S�B�\`n:�c�F�c+�jB�0�`�r�PҽS�X,�0X �Y���ʍ�}
�B��P�0b� �� ��Xz.��e�,=��D�0"CK���(\X.Y.<
����EE�=���,5�5�M��e�+����)�S�����ʴ,PO��M�J6��
]a؈�4�J�a�`XEEঠU���V z0��`�ܟ�4O?�N�t���BS�\X�AS�\x��}��8�Xq`"�cb�9���*$���_��S�T�,��弱�f!=��
�[Lh�^h�}^����,�@x�6k��v�����(\X.Y.<
����EE��.x㠗ā/��_�$�I�^�a<�~�@a<�^Y��0�KYz�	���8�s�U$p |u�@ϥ/�@ϥWp ��ҿ.�@ϥWp ��r(������<����n�>�j����Ma˩��ui������6�����'Q3c�#jfL7)G͌��P3c:jfL���fF�Q3c���Q
�4�tV������O`?��H�{���=�Ӄ��h�)φ�,Ee˘�C�����m�>�������73�����QS�*�A�����IO16�
Ά����	L;p=I�uښ��!���G���Eٕ��u2:��>[�xV�k�x�)#^ d� �@�@�x��$^ dV� �\�2�<��H5�`3�'3���� ��?� �P�`���\#)m$x��{¢kd�g�F�|V�k��O��p��9��:��<:��t��Y5~	��u�_E{��5��'3F�\�g��.7��c����������ͬĶF��d�dDv4.;�]���N�e'�Sq��Sv��̫��n���O�&��Dj�Ô�ȩ.��P�\ڀ)$�u�}p�&L�m�@u��o�m�a���Up/'l��M��u(*����0�8r�;�2`��-����~��
îh�\��b0��P�t������7���1�b�I��ҁ{H[�p	M�t_ƣ=�Y�S	��s	��_9��������>���W��Gd�4�SO�,�,�)45��7* �m?�� �n�.�X��[�3�hf�] Q�� H=� ��b6[�,���d���RZ���arOL���*1)$&_�$��L��a�4LP�	*0q���<����$&n�d#�Z��"?��l>̈́PߠE��Fϸ/��[Oc*�w�p����'�c����X��8\��i^��p���4<}���a(L�z^����M�����[?.���_x��!�!r:DwC�t�������!���Cj7�N��nH����"7��ƚ����Ӽ��̗��]��r:���n��"Y�p��Z;ۖ(ͤ�t�(Jn��T�)��\o�4�t��~�L���V�&����Aֵ�ά�;��9��^��z=�>�߾X�f�揑�M�D)�y��HʱTt"2F�t=h^��>˂�4�M�3R%S6��&����ʒ�»4om��P�7-��l%m�ݩbVs����	!r�ǚ����I���!=:����Ѓ��!���C�����R�!I�CYxHn�k���Tp�/�f��1[��ޔ��/�fD&�9�w�j��~���pq��u=[�w��0���>���F�)�,f�#���n����ώ��2�u�+[�2[��}<W�nf�u�Z;-q8�`���Mm�s������4U���_�Z����T-��RN2%2Mv+-Ɗ�IF2��~�����}�r��y�d�1�n��G��/PM�_N�C$��!u�l�#B��N��eX�Ѯfۻ8شr����iD�-�d�]w�������@{G��g�f��Aұv^�hMy&�Tk�=��˹��9����^�=�^$��_�{�����1�ͩtB��4G����o{�~�y�N0���Cn���/͢\���M{ 呐�ؙ6���h&:ݚ����YS.���P"�2����Ve�����-@*k �o�v���[~	$�oSOT�xFw�'t��d��H�عIv�T�\�e��J�L2�D���U��85��k *�׀g�=g��o��n�Wݎ��f�a���È�Ǳ�| )=�f?B��k�ܱ��o߿I��+�./�)��Dw)4��J���̅d"��G��h))I�����~�J�*�����MH{����s����������H���,u�x�����G=��J�ST���X��0��UI��u{ʙ�ʔTR�q z�0"��@z#��MǕ ��Kɓ_�����`񰼊�5�2.뗆�	�3���q�KU)s�h^��ڰ =6��̓K=�,K��l�jv����;;�;u�������NI)��0"!��Dp��v�m��c{y<8Y+���Dp��8��i���ch��c$2m��Z���x~3ڎ��p?ЇY_�[n�{�VhĘ�PE�2xS �%L��Wh/�Y��s'���͹;ۨ�;)�1��̿��������0ŝ-_>V��v��������7������T������Kз��r�^��-^������fvQ�e{<ڰ�ͧ�b����%�t���b�Ƭ�^�oooG����z�~j<�ʟ�y����J>bj�u�?�b�%�2IdG%��w_nG_��X�@dpH(8H�GS�����"2 #=d���"*8dp8Э��%dA�!�Z����!"��G���,��>D^Y<p���Ȣ��G��%a�����,28XTpd1��(hׁdA�!�Z����"��F��,��>D^$8hdp���Q��`�$a�����1l3�]� �S�9�KȂ�C���@���_

��a����QB%��D��WP��� 1@�X�~�� ,=�M�.*�i���P�g,ʌm����A�6un���-c $Bc�'cz
�qI�0BG}\rQq��� �A�I�* C^D�嗀 �k{�lˀ�� �bٖ���G��D��$��Ӧ���ʰm��] �WoW�1"z���}�����0'���N_�l�OB��h�iyXQ7v�Mjx@�W��{er�။�� �q\��5T�M�QUJ�m�=�j�xB��g�D����k���r����p�`<4��)U`�^]`�y�q\	���HUeyJ�1�+-��y2�-�×�J�ͫ���
��Ќ^@�u'A���i�+~��dNDh�?�E��eV�C6�e�T���;�iY����#��b�������������Rqx��M	%F�QTQ!k`�}�*6�����A(�8����wS�b����1VڨЀ���>�����h�hm:�JwW���8��FAU���Ѐ5�þ�����!����Պ6�T�� �C���`���]�puHw2\�h��E���E�5�U��Qu�����>��y������fm뙙�F7-��`�/[~o3���jm?����2��_PK   �beT��/J|�  v�  /   images/265b7ddb-a887-4736-b161-f7ff4501cdab.pngl{uP[O�o����6w
w��h�"ť�((V�w(^��ww-��^�����̻3wg���=��;g��U�C)�  ౢJ  ��{����+y�����NA�  t��.Z>�  E���g�^�v4��;��"/�������Aَy�u��;O|+�؆ױ��`Ü��-.X&�5B
��]#���I�Y� ��`�v���y~�����o;%����/�/��^`"�#0��%��s�i4$+�C��{��b�>!���$����Z^%[�%E��\���YM�  ��u�c@wVՂ{2 x�[���ٍ��ۺm_�ˈ�b������C+��^�L�-і�]���ug� u�;�Hܢ�'�xvLH4�$ �h�~�D��H0}��ў����z�.E9^l�<�3�̋%ԕl6�l�5�b�Fu*�����g1�1�(g�?/bi-R�  �꙱J�)�C8i|���E�c>�����!�~�X��>8ZY�^���~`��=�"�{�<T�����)gm�R&�����l"�"� fn� �SH�;T����0OtY��}�R]޼��Z6ړ�V�:(R���R&�F�42�/"RP�����t���G��x �;�"�-�<ƺ��^��N�zF6�BԉÐ#�a�D�f&[��h�D2�wf�̈́Q����<�~O��q����vd�h^Gc�N��I�`��u0�QQ���>_w� �ٺPY�>R�kR��艥��r����?�ԡS�D�?�y�~��<�F��\E,4 B�����<	�����/����0��u1�m�?2 
F���C�F��w=�t����d�g�赃@._�Gf �\�n�^r.��Ut�� L24�^b.�X��ޤG���_J@���P�:�����d�&I̹b/��9����we7Y�A�-�S�������V
Ǿ���܇@ڍNr��3U�'z~������ݴ	.�|�$F���+�^��z�$`�@般)],�]"�ō������2 "�������v䰽g�vw��z$/W�鉸���,�EF���=q������]lEv��͎��1���D�w����.g�4��/�,k�c��}H&e��I����b�N1O[�������x+�o�)
��,�Nr�rYbu�����[���?�n��� �i8�����?8��
5«o	��vR����9`�У�[��m���թ��99pH�li:��u_TQ��lE<����~ܥ���H�@ɢy�H��þ�h��R]]�p�$.�6P�/�쀫0s���Q��� 7Ko:�/�Vi��XZ�� 8Àb���Z2x٧�>5����>��W��o;1v@�N�`��T�) �����耔��
 �x�'�G� �S�ě**�D2<ǚ�_j����meP�O��2}!N�:!�jώ�3d�����hk��X\������զi�Ŵ;�
�.�36S\t~�_=s�f~ �y�c�U1[xs�d�&�t�]��t�G���N<I���n~a5��1�-��&�	����.���M�iz�Ƨ�X��Y���;�L�LY���0�G�[���\Ƥ1�j�aG���n��gh� ܟ&�#�o���x�������f��?E6��{�� ��G��Eʉ�r3ͽ�Zp�+�|����сK�Ty���O��E�M���B%��-9<�������������xb?�4�R̺���r���ټ��E��@W]3���n,�,|ګJ�;���Ǟ/����i3�����z\6�����f�����t�;�o��E�����H2��+Z�k�z�j�6��p1g&+�����I�h��,���c]V���F�>�����$f�L+^�=���?���6����ZF��E�5?(�o��>3�J�%����qaF{�D��i�Ծ��8u-T>��Q1Ĩ.�f��QD#���7�ɽf�A�{�q��]Րn��xc�[�ǤS� ��S'��r�E&KN����	�DE/{ӤϽZ�.��=E�I���kZN����
�%?���L��`���;4#橖�bKW��M��}��uh�\1�n)�M~a���otQ��4�ϑ]RK>,��W�md�8�������[=��i��$�Bh����DL�� ���#i�o��j��k�V�����&XA��r���.��2ف�/�n/=1���v������C&>��s:q6ԋo�3ۛ��0(�3W�Y;� �+,���m*���p`��5(�a�Zv\�b=��]B�ڿ�'8�p8���΍X�M#v���3t���#���'�{�pyX��?!G�$�]��W�!������:�|g��F���S���opP1��#~m4����%&����h� 7���sה��3��D֗E��ߟ'L��݄Hj�Ӈsn �I6��Wy�BW�B�%wA��!��~$�e�X%*&�`�= ��X�	�� W׌�?cT���(�-9Z�'�=����\ћ7ݹ�f�^�n�#.���Χ��Jm^��
�>��fGJ1�������?+1�=���8���Ep?�B�s�R�æָ46�{Sj�5�;�%�KH��a�������ˌ������"����4�vm�Qe	N�%�__�H��KE�p�*R�c`P=Z��\�!�����Dw<'a�$;�L�9�K�,:�Z���b"Ƨ��]ֽ+��W� G���!�(��;����a�m�ڼ�=�`C���Y��9��� ���&��8M"WdSMy�w	��*q��wuǛ��O��j��7g��L�d��p�9=	*s" PȧLL�E�-��Z}E��X��y����v:L�j�@i�:�ii_��R��oZ�w��w��\����T�����ݱF��ڤ�(����듼�tK��T"�^4�-'���N��=vb�*���-�{�}�'0a1 �^/� Ԭ�Q�`���(���9��Ѭ��$�O��Ĩ�D;b��Ö�5�y
�ɑoqT�G�qQr�����H������Ƅ���|`?���f�E��>�)r�K"�����"��6�ϋ�[����q���V.�@�u��v̊/j�^5�~�(���<u_`�Be��L�7Ff����|�p���K�n����w�wq��j�}�s�^�]��TDA���9�t���(���>]/�F�{�4(n��e�����0��̻�`�%f47\.�cǔ����7}�]ŦҦ$:5hʯݧ^)Jܠ��^��JV�C>]O�L��� @���ME�z�/��I�2��7GM�z�oKBx�9�����������Ӓf�I�@���1��A�����b����7G����twS�U��z��Yl�6#�ͧ/�֫���tjM��|L�id[�_]E�o���tl�1mm�<��!
�	g��n
��� �}��S���M��k�?h���G7���nwi����E/u�q�Kle��ԛ砸5}(�x:�0�
z�`d�]�l>�L��@�f� ���|���E�W�R0ز��mI�WIb��4��s�φPpP��y���=GV��=�_-]���P���9}�w�9�k��J���ˡrU���	`!��{�B.P����K�&N�"���E,"*%{%R[+r��d~޷0(�QY�9���An�9��a�۩����;g�����(�.9_v���!! Rŝ���n�{�+1���@<�qLK�ܵcU��n[���,C7b}YO�G�w��ݕ���P��O�� �ƞ:n4��|�$���mث*+Z�/����i�D��-�
��,37V'�;�{qQȌD�w��EG�{�㣕� ��rRl�v�X���F���#��uJ���
��ﰈ��hS&��yz?oC"H�G��tiʏD$.$�Eթ��2�Ï�����-���p|�Y�޲����� �����d+�����o`(���>Q�g$�O�je&��x��Z�}����H	�ڂ�s7�D�C1�İ���?��mـIz���Gi�-x� �N��t���u�ثn����MS,��Ј��0#�o&Y����SI�>������V�`�%) �ۇ�OZ����+��
#	�×���p�hHQa@�x����a��zv�f�(�J,i�{?����u���'�@���PU$.���^����i\Ώv��'�A)����6{g�OORX�^}���@�|��ZK߫�����#"�n��c&w�n���1H���9-�����/��J������z��{<��Ϣ^�F�b��ڋ>�j���ZJ婐h溑˙�@H:���R�^;�skm��� 9*���!��Q�0=ԗ�Q��T�B��"�ψ[6�"	K�c���Le_�N=a�^\�Khϗ�l-��KX��6S�q8K#]�_H;*E�ABV��H��K/����x=_�*įl_p�����M�0�{"2�?��d�����;�VG׋n;�����K�%�Q�V[���5|Y6���α�kK������9|=��zD�iBp�R$iN���p���b���[g�N�(�J(7��k��Li��]�"B� �i�:�,(��ˢF��T�?�8o��褫҇�T)�q���:�[��[��C3@���5f�xğu�5K�����_�q�(�����.S3���FO1�0<Y-:*��ktI�W��|���0;��m��vV�����(�y���.�V���n�
��(8K�k��u��:i��m�")ճ�(�0��ꍾ��&��ĩIGbx  � mX�A�3{f/�M����Vb⟇kh��e�sk`��z��3VS��/t&�AB8��#-W�&)e*�y��0nZ�ˤ
�N;[,����N��ڪ�0�r��٠-u,�Nޮh���O�qZ�r�/Eپ���m&���+��7�K8߶Ϸ-����+&� ��w�pe����"����O�V��8Z������1lu��$��ͣ���5奡� f�^\2�?�hv=Ya��<���Vd��������)�s, T���|̥bZv�~�ng&�&
�Ė#��"0����|A@-s�Д$��G��?�P"'�?mJ�T�������3�Yt�~K���I9���� �G��63=��/��4�Bb��JT�z�T�c�Q�C��SZ�@��l<�����m}��`��x����\��0c޸14��2@�m.U�+�Y�U�yXN�7V�:����'���8�Ӎ��3�Ħ�s�}CŪ�0ӯ^��PW�f��!�C!r5��Z�B�E�C�瞇P�(��\ΉN�Q���~,��&
)���bI���ӱ�62="����':��[�M/[$�Z�
�H�YHGc��/���n8 ׸Q�E��x�+��x��u��۠�|�|��@PH�-j�qC�g�-YҲ�qC��>>v*��z�N���l�!��zv}=���3���x�%���K��o5���Cbw�s''�>�����g~fk��0)@FF��?I�	��8.����*)�����B���b��^%2"��s�ƙ<6�Sȭs�g�������YP��j1u2�LNI���x9�@���kN�+��'�t�%K�.���`�2�'��2����
�LM�SA3sh�T��)�hB��:��J�ye�@Ir9( k�f�nm��W�=��f�䓴��4T��  ���J8���7q&�s���K�T1�B�� d�!`��4���	BY+��O�TB��/�o�^�a�[i�[�N���@|B�Y.á����o��z��f�7\���ҡ��Hf�O�ᭉ����@��k��Q�ʥ�s�����Uϒ��'���I��L�& ���ӂ��Z��Z���2�"�}>�e��'�b�Z�7|2�	�9���@p U��'gj,�9]��-��?\�K��AB6ն��@&�N��]�͌ۃ�$����ݳNo?(�o��f.��C��եXܑ����Yql|B����f$"2XJCB�r�uх�ˠ8һI�b�~�h�<����=���F�wœ\n�ν�!�Dޙڥo������in?�PMUE�S�;�<ů�m�U ��T�C~y53*�U"p7��#&qƷ�x���;�':�f�fw�����JT��d���%W�%&I+�r~��I�1DC»���aQ
�	��<"���N��
���Q�k��D�Tm�&2lw���͕�M3�a�)U�����{�C����{=ccDZ�g!*U�r2�S��_��&T�j8?2��y�
�k�P׈	77�Z�(a+��	������[��cǅ��K�&v��x4O(9-�*l�Jy�ąx_�1$��s��3���E|�r@��i=󛵫�J5��s�6Ɖ,�`]v�qDD	J���T%���%�,�>�`�ڄmM���{3�*w��R�ѐb������!�����A���	������~�\�p6V�9��D1�ӭ#�F7��գ����UD��V���/J��n}M?�l4"_Ekɫ��=�U;�tu���}���ڃ�2�T<4�U�'t#�}�u�U�$��1���~ �l4 <�%�#��7��&���wmD�[�#ڸ	a\ző9�8op{QR�����ܺ�b�e�
[-8e�b&���M��:_i�V�k�7�?!;��aQ��`��L8�bC$��I����Y�O��J��W���Y�����]�)��y��@��f����̌~����B�u��������_΂��&E�ߑE#1}�����+��;q!q#+r�Hi�|�@Ĥz�%/q�6�T`�tz�\L��+�|�m5�2@���?��+���t}Ӥ�u۬a���ts�;�R�):�sc4o�IMwU���4P��|�2%�4b��ad�+��0��?��ҏe/+M�W�X�.>�US��wnC�����e�K��;�!��;a� A��-�
�o�p��a�ق����,�*�U"80��F�e#����S 	�f�*G�m�`G�P|�Xl��>���ʤ ��Mg�X��N��Vt�^���q���g�#�k�3��*�2"�;��u,
L|Ϗ�Z�w�W������k�
�22Ҿ>v;]	}VRV�0�o8$v�gW�x}��F᠓����[��.�q��'ygܣ��΢T��J�e�R����aQ�zB�g!����*����0�с������ɟԌ��K��y��nl��IhE~�-��ᅫ������8���N�K��b�WqS=��Y����z�f��c�������+��ޕ�`���W�0��ޮo:~�t�?	}\��&����V����V>����<��f	��+�C�㷞�Xy�@����V&��YB(��^�>�Ӑ#�Γ"�������Qi�gI�VFy=�t?�N�R��&@r'iYp0�wV����_ͼϜ����'���)��oʴ������(5�7M�|#�������+��%m���h��9$zTS��,,qr�\h�lA�j~��Ǒ��%�v������xݙ�;�)����O�9S��_ɢ�����뛳r���OC���������ȁ�85q���>������sN�U�l���d-�&�	���7L��7�>6��'{U�\�n���׶
j{�?RV��(�
��R�rZJm8#h�*u2�Y�1?,9>iM��tQ���O��Wz���>"��?J�4�,�v��}��dd�D��*�2_�I���_9���s���q�8�'Swub�P��p�ID%�����i�L�4�����{6io�x�_u�.����I3�LQ���� ��@k����Gч����{�ɯnP|�c�.ʯ_��Іg>N�k�3�͹uFr�,��*!6���g�7��~P�ΰ��a�p9~�m�YZ�]�){��o�W
�tQft��������ܩ�{�wqH��#���bP�P�`���(���ɸ�����=�x��mSM��������r���F��#�1�|�����+U|�CV����@�ce.����W���N��3'B3>�{��e<�?�f���Z9Vj5$z6�t��3t��p#_�Ҭ���f;l~�q��u�qxw~8�<�tr."�4t�c)`��&ǁ�g�������o����k��UL�U�Z���|�.E��oxƅ�S����滜��?C��3ւď��[�&�|��Z�2����6\�j���34���wvv.�O?����>���T5'���]�1gn#�̉�P���2���������d!�qA8������UV6׶ �fPc����Ƌ����J�g��x��SH���0П`E�F���dY˂�{j�j��'Y'OYn�E��A  P;X��75\�<�'4k]>��rj<�˰�,�Uǥ]9�����l�op��dM)�Ɠg�1�}��H�����#���d����|:AM�k�˩܉/�����t�չȉ���Y�D�V�� �H�|��l����ک^)�Ǧ�����伡����f��YGY���:�!��:;7a��e�=,.�K�E���n�ZAA�PF�;O��J��˝��)	���+�A55�Z���;WK����z�����Ŗ�Y6���8�(yV#~8�cI�RZF��zU�Osy��$���y.�s/���}��d:O�����۶����'�sY��k�#����ac�l)��L,�lt����lF���r���gFM��:}5��v9PB`�q)�`ʐ/؍���ѯؒKwlf�
��L-zޔvL0D�Ĥ�]��[���c�/H�]��[X_�|�J���k��Qߐ����s�*]�lЯ��n��ߩ��'|+/-������sk��yE<V��	�	2�Pd�G��d�,]N
�841
_����tY�ƴ�}�C�Z%��� Ɋ���k���ûż������2��q�ퟕ䙡$҃�檺�f�a�����OKM��	k�b<sf�oQOgK�&�ag�ķ�r(���Wީ$�o�.?��{*,ܩ��)�4���~zt�{l��D:���"�8a{&9���.�D�ym+����҇���E2@^��9N,s��!�䳹@��������߂��e;�53��br�m�)W�a�f&��<��?ݠr�pʡ�~wh���/��wh<_�"�-�,��K�4Ф��ц��zn���� B�bD%���jէ� !u��
��*�1X��8��34.�$���a��k��Dڒ�})�R`YPz���ݫJ���QQ7}:=d�W�9����v��t�WU�q�I���\tB���<噉��_��W�@���`OOK~;&w�du���t���DB�Oߧ�+�4r'S�_n�צZ�7�O���-�t���J@)6&(2>�'�U�.C�G�$J�8y+;�8������N�_�*��z�*��)cvU_��R�j]�E�R,C�+�,n"�8�� �s�[-*"�b�ɠ��<B�}v-7������X��	~p������ݔȐ����A�D�_O���ۚ�K}�l8�$�O�h�_�ؐS��Z��e���3_���s������q��9ĩh 6�s���S�PE�ҍ��S̩,]�t�C`M�3E���}�.�y I��4����D�B�J��1	�h/S���6_�'LV�j�B��k��|�/HuI��d�I>��;{��p.Be�k`GLN����Ra�A��"�)JZ�XZ���4�b�)-04�^��m�,�Z,�B=�ʞ۩E��O+Uw+SL��zns���k�������g�������3KWKW�-���>��A��r�_���!��MP6	�T�ԯ��*h9 �a�_Ck*�;2FNOP{AX�?ڎ��P\^����Zioo�5���+o>_�?\�ћU0`��[�����ʧ�љ�i>x0!I��p^�[Ґ&�})���Vg�β����T�1��Y�o��q4C��f��(Qy������TY�R��-��_�͚~56�D-��C]\8�^"��o����Q���p=8�v�7���~sT�����BJ�Gyi�F��Ҵ�#cl�cI�فZ��4G�W̡��������rz�w� �ł*��2��V�ʆa�W���\��2��w";t5G>�N�3����j�#���;P�h"Lf�#�kE���9H�������yo�I��}�E}}c�ܢ^��Qb�Pc��	�~H�L���R�@0G?�R3�H��֎f�8�^�.v�Uʅ������"=���&�`k�-w��:K>w��tu����Ľ6���?���TW�ہdM������VOj7�W�<�3nfBM�}��>��9��u95%�U4w(5(�s����q�p�n���ŋ�����[��Ek���������K:�]���?,vt "q��5%�ˡP̤���沷��;e��f������M���e���ǡ�zd�$��Tuz����K������[щd��qD��s���#������Y�ۆS7#���K㸂��x��bi�� ����{��6��D��~X�0�pygz�K|
�zM�(T��+C��U�6�݊���ֶ���?�/�&���Р�2t&m�݋���;Z� �Ҥ�p�l����l�l/���h -�E�/[���FBM�m=����g�k�Q��VԶ�������	�E�r��������O�q�Tn U��x>�*�����{SgӜWd���S��ݬ�גyM����2R�D}6���^������h~o�l��+�`�gc[���'���c򀜹}����?�i,�u�f�7��_�����D�m��L;%�Ir������b>
��s�}���v�^�S�	^C��WIy����m^��2����3.�j���A���82��)�ٌ�v���}s��?<�<^v�FČ�ܱ�Hi��{X7�P{}�.u0Z�]�8�9=�65��~��$G7��񍵙���^�h��+�����Z�ZN"b�ŀ����	$ϡ91��ai��ɞ]h(�h
��W��|�I�՗��qf�E<B	�[��,���|�s>==b�w;�f���^�Rd�|X�(o���㕷T��0��E���oϪC����lM�T�~v�ro�����9��ٵ˾�F��Kg���U�P�$]]������?�Kz�S��{��®�,sT2Z�5�����=섞(?"�&���MB]�=���M��n��|���� �t�YB�ل\bPe��6��noW�f69����xI����@�I��^���S�?��O9.Z�L�����4%���о��3�č-��֔e������k{�_�>�-N0pxa����h��"^^�K��z��+Q��WS��%� jh��Y�B���ɻ�qNy�,BT����F�V�rצO$̆�X��a\O۳���k7tH;�O*�,�⋀-�F-���njM���,�f�)��vOj�3�����y�y��N�X����M9-5�,��;P<���6_�ߌ\��pu��J5�w'�j��q��X����c�Ʊi���,x�x�S���&�%���;��5�����Y�����q�^�7��Y��ۿ��D����@��O�����Ƚ5{	��H���mߑ��$��j�� ءzX�}p�T����X�rp*����X���yv�w�s!(MZ3?������>O���;�_���g���h��r��~�i�ʑx��Jڵ�9'��S�x���� <F��)�����车���e�a�3%Č���vx����O�4�t��U��/@$ԘUj��oREۮ+��Y�GcEue�F؟�d}��ל���|�J���O��b�hjP����/���W�������r�����ԯ���\�����fɄ�,u��}���1�]��;�������2A�v#�q]�I���X�÷j�Ȓ���䴯��[#t�q�M�K�����TŻv��vL�����/_>z9�����9�����v�AYY�,78���#Ҧ�D��TR�@���Y7Q)C�T]Y�y?�}P�N����8U�"T�eT�]������*��E[��݌���/��5#�Ĳ	��"���� �:Bz=��J;�܏��ϭ����f{b!�z��dn��Hഭ��;'�<&�t�J^����ܡ���	l�#p:'�"@��a��?ha��^���(Uuc`�2� ���-�Q��7�� �)[��s��,@��A���t�::�'�������@�HI�GÕJU�%���UVo��PP�T�'-��oT�դNK_u��b]8�JNt�w�+B���۲pͫj�Մ����V���$Z�}�ÖΡ���U��܊T�����A���J���FZ�M6]�Y\���xe�)��݊�/��y����{�����R߮F�@��f�� Iᆥ�(1q��+k�Q$��c.u}�k���/��|N����.%���w�k<�a�"�P�W�;��e�Ī���%B!P�@d��4�(��fN8���[&I�Ek���u�
&����W�T*�hȣ�N[)IU���oc�G�EB�7=O���d=E�?P�B*�G�衯7����qH��hr����-��J)12O�9L�q:�Zm�a]z�0�&Ri�˔�:j{*
����1Tf���d������U�8��|3ɔdooK�˞���ؒh#�-�axxa�$�piuTP��|��&��ӳ����j���(D|��
P����Z�����̓ ���U-���O?�KL�g�"$U�e��ﲓ�H�Ax`
p��v��Tb)հ�G"/.�"-��%����p>o�I�\�z&�1L��x��È� ���t�(e�%�A�+� 7�x$��TV�2���Qm�I%�y���mMaWQ��M��
C���{]En��O`����}`���/b������m�P��X�CҎ�@n������;�?Ds��d%b�^f�y��?p@�(py��҃
᫤�}:M%McKc�Fj��,Z���Ń�)�4�#��HѺߪ��~T(�`$��$K�=>�4
��2���T��L)����pxjm�أPbV��0�����h���A�I����JoLM	�3=��+�yn�tN���8�ǰv�� bZd�����/8K���j`1d�EB�:|�%ͪ���TӚ�4��f3��M._�Y�Ar����q��%��4�h�V;�tӽ�{�֎�ܜ���YJ��-��`�� sr��i���M��� rYah�FV�}�Cl>�,ܡ0��gdi���s�G$�`qП��2j6d�hn���e�Sbݑ�H��n�����t62��}(.M��o�8B�O�bZ�i�L¢	�d�~��
�!����Sڣ�Y(pb�'�g����Q	�k�����m��m�$⩀�9�u^o��)J�`�|����'咆b��m�]���'Q�W/�'^��[[��Eˀ[����(P*��^,�aP�`4e��S�Z_�	gy�Lh)U�aeB���(��ܔSn���/��F�فM���nt���0{��R3��]	!����oǥ&N
�fٌ������盔|��  ��hx�y,����Ƶ�S6�#�����
�A!' n�?�!�,�0� esJ�	0���0��O��eo�"-@��Z��[��!�!��'���gc.}%����~V`$$��d_{�c��K�������Y�)�6��H��y�{I�.���#��K?E�!�+B��p�ۿ,;M�)��& -n���%!�n��<���CE�0��|��1���G�P,����"C����)��I�"B��A�0u������8�+���C㣘��<rA_�:��7��gIV���E`��R)��%��cA�
��dX�Ez/4>;��-g F�--m��,j�Ӓ�?�l��$4�!0h0~�^��>��/�X9j����jK��-��r����ʨ��?Hkt����u��B�CX���Vd�<�y���8gfS4��Hv�@���1��E,:ۜj��R���$	���4ĎpS!Á��>�@w÷1\�p$k�4V��y�S�_iI�_��\���#��0�B}�y�5Р��p4,��Άx���q��@�B���#	����/�rp]��df�c(f..�Y7ET�O������a1�_�wi@Ș$�jp�x�7�5x�.��VY���դrE	H�s�3`�?ß I��1���Bp���
 ��Z0@X ���(�}Y���5��/(2#c���ezeJA>@��Ш����,��/��ߺ�B�� @!	مLf��a*�{�� N�xីsU�0����6=��� �g����X&��ihf�_" �2ʽ�ط��i��~@�閱u[�4N�e����.*6����ם(���t��� �oe�_\��Eڊ{z?'O��^K�t m�q��(e���^��\8Q%b �-؊�zb�.x��b!��(8~O+օź.9�<�����ӣ~�"I8�h��C�)Z����5� �����e�)@�F��fp��Rl2|�p�wڪz���:��K��	���̳�Z^��w�������!<%��o��O,]���u�7b���|���)~�����i%��O⯀z���.��J�_�[�o��)I������3����Q�S��U\�����������V3��f��3L��f�y�=t����~�=<��'=f��n_�����МS�do';L������S
xƙ��f�V�H=(S]W��_ב��z���S����#j�������������y����T70�_�tӸ>�Y��z����ie/N�`?�gI���t�?����;��h�3+u���3Mb��럴i&n��7�n��>�@h�����Ō���i?+����̕��������m��̮b�LPuhs����1Rz�%�����k�{�6���ӻ�lc�e���޹k�#ZO�^��B�L�rV:��IB~�h/��o�7�e�ܗ��\�Ҏ/rc<���,b͐	&�A��Z���(햡:��Q,��hA|������0�e�ѱ�#-�)m5�	Gm�5��<�} ���\0�<��싚������Q44{j
��1���߈Z�q�v�\v�����)�)��(5�~�)��q.���Gm����
V��p�� �Ľ��.VeU @�����Jvst��I������@�����R�^���ws-�R7��ϔ�{>7P��\)��{yc=z5Rz���-�n��xI}��t�A��u{��y�)t+�_u^4��VG3�K�\�&Pt�r�}p|��J	,C��S�$�O�M�Z�����X$����辝�����<I6@�,Q�A{¸:^o��|A ����s�ڟ�nJ[t}��{�?_������C��=�N����s� ��i4>�2y�/v��W�^A߼�h�E��oz��	��J�:�#(���,���PEi��E��c��<m�:�f���(��'��P���] �Dc@h�)�)}�;��Bѝ�ɟ
����
�nu��{�{��}6��U��b�)_�e�i��{���7��J����9��u
�Nr����tF��fT{v�@xBe'<��8���KVKjw��N�x��n�O�Ӻ8�Ƶ��/j�Ǜ��s�Y�[��.�۪ �8,�fL����و���Z��VfW)y��f_��+�tc�'�������@��h� Q< `��BÓ�;��V�g�0�����TZX����3��l�s�-��XZ�6Ţ!ƀ�LI@a�l�� ��E�
���m|�1�R�����#>=���0 �����F���S�iI��l-"f��"I'��[���G-�0�~��h��| ���57��Pi�]-3P�b�Ux��ժ�,��f�b��1���
l�>1o��,1<�zd�r�/�23F�̙!W�%��E�)�2	GL�Uf�ԩ�.T�Cv��`Z�45��Ǎ�(b (&��j��F������nN�C�ݤTvu���$�swY�i�gp����*]h	�'�L@��GK�P��V H(�����4|�� p��X�π�x�d��a�R5r��#���u�:!d�J��ţ�Fqw�:=4�t�����q@�r�c֑�~'����U�%EPIP!�ZH0(�s[�ez$�s6��5(~P���@�HQ/r�� �0m�C���u���hB�M�	'�S�숉̽\�\�J\��z�p�Y_z%�'�R�.���`>7�%)QT=	��`�+{'�7T�ש�7�'���С,�T8l U��������T��N�B\���B����: �9	��.2bc�p�(�3T���9�^s���ƕ�i4Yr�����X�@6�'b�;�/�<_���ըA84���8Z㢔ۨ1ָ1~��z�`���}x	��.�轅h��`�%�j�{��ktщ�Cl�,�K�X���^��^>3ߙ�gg��}����\�uֽ���tb�S����_qk�������S�fg7F�.���7A�P]sΣ�O���v� �j����K��7��OTr������D?�G0m�FagDF�Ͷ�Q(dW04c��b��5`�r�U��0Y�K1��"��U��K'�� ��Zr��2+�R,B�oCB��ؘ�I(0�&��ɭR�;���5���WЇNt���� F�t����q���_۴���Ԣ)��GW�Gˁw�(��4'14S�2�w<KSw����ل(?�ț7�M�^��e�������>o0ИƇa��XK���G��Q#<�k��@��qj�ǅ'KB�� '�8Ħ�e�*�_����A�Fԃ:`�1��IF J���;l�A�7X5v�$a[�:��ω�CD�~xm%��Չ���<�ɸE+���A���4�`tlLlf�IK�J��}*�N*L�BOrZb��������CeYB[eN�b]	L���B��fX؃�/�/hK�9-�!�t"E16�;����-�����ضPE����0_�f��G���U/m
����@���hxDh�ĉ)22/5��CT�NN���L���~�%UB�"'o�����#a`�W�~!pG�� ��EI$�jt�2a��3���1Y�]1a�u�<3Ta;��mk9\��>�ד4bZ��h����ɪ�ص�C�1�	�"�0S��;?I�<0��1q����e$��rr��G����Yv��3Al�~��e�2t��x컷8.���a8��v3E����8"2͖����������/Tե/�Z|��i^�e�4J�H�n�?h�:j�<?�����)�>�$K���J5�!#���_e��f�J9,[Ο�13��Ph���ؤ��3r���=e~m��a��0��&�����{�|`&4���(���{�4N+zl��r+G5��"}atpu،��g�޲*��}�vvT2�m��u̵�49�e�RB��Hu�9t����LB����Wm����Qk��!#?��գ�� ei�gj`v�ĉ5y,<G*�SU��9U��f�|,(5����4��D�,��m��I_v�Л�+�G�G���AF}{�1���,r�5�6���D/��Q��r	��|���gRЂ�e��#���8�����T���F
�M�<pF�ǚ/�F��Z+=|ɞI���JC��UOJ�(�!���5�h�|� b/R��$T�3��jVMG��R��>*��C�2!yP�C�L�Yʓ���HA{�NӁ�T���N�Թ���/qxn	X]�Cq@x��5��P��<�Cʯ�>тڕ?S��/�:(�:�7�X�~�`.[��tO�/�HC���KB��<��~����=�H�N��l}y�lǔS�,��?8�3�(�Jr��7�]�`D�-�mk�n�q��]��6NL	P��K��W�c�D���nFAU@�pjF{͊e��I�3�4��K?�j����(a2k��Η�0?��[���'��P��\����4b8.��1��R���P�H����;#��5���[-�ZȌ�)1�
���$Q�ޫ��6U)���"	�R#��z��ƭg�a��q[s=�w���Y.aD֐UzZL�k�b���x�p??�0m]O��/F�w<���G�K��o#�`1g��B�h d|�UYY����`��)�_���]3��H�o`��\���\�^}���6O^�G�u�ѩ��*K�۔��n%��ѱ��2}�$.�,NqӨV�Y�2X���
��e=-�����|������V��O�颛����=����?�ب�;[�i��'DN�;�It��=Q�7rY���Q�=���%N׆Bti{E�pЀ�ͼ���ͤUa����M>G�P`������I���q�D:��7���?0>{��leL��v�N���5��bq�?��D�`�'�E��7��ck�r��v�CCW�}֙��G�ğ�����}����W�jz�#�A�>�}�jk?�W{՞#�Q3���n}Ǉ,_+)]�̒�r��~��S,S�ٰ�7T���fs��}�N��PQ��5j���E1�������������3�u�f�od#�ǉF|�7�k�hpp������%����֯���P�2�U�8r>���]�W�8���-YY�M�tIn77y���m��&Q�Ç�l�F��:��*���z�3Pd��NQ���okF�=���"f������/3��:��b������Xs�-��/��?�X�m��>�}�T�Y�V�k/��� x��8�z���o%p���4[�|,���<��t��sI��(��C�9�>/WW�����3[�F�~�gY?�ؾ�XTT���i�MV��|7|7/�p{{}Z��y��	q-�[����4tB���Uja�ˤ�o���z��!J5���K�`��o��m�£Q^�IVX/qB��a���'�ǵ��e����F������7��^�}�3eP U�=%﫭����s
Ndw����P_�G!~�PG �jX���n����V���W�T�@��"�m}+��I�="%���޳����%�n8�n��s��}DǤ��e3,�!��n�s953�������������Ӑ���=-�J�Ֆa�2N���6�f���_�2HQ�=C�;�Z��(��o�g��
��������ޚjq�c3,����srfmr;��}������;-�w����=��m�M_Z�6	ge��������U)qn�Mr_�/�}�p,�i%&��[�`��l1,S4}��U�[S��`-eJ�c����v��e̮�'!�+�֢��h��P�������k��"#�O��h���n��er=#�۸��ɟ6�"s@�����.mW��V_����ξ��lo��ka�ZU�����=���ݷ��m��`����K��Dlq�j���%%��|[�������'|��+R�=����'[��ڳ��V}�m�����F�;����Oi�R�(X&$T�r��JEsC	i/}!.� 9lB)ʞ2��@#[��J�R��V�Qp�yz_�����'*���`3c��v���A9=�������x
)O@,���s��o���{�E�R��Ka`��O�w2ȅ�?P�oswrǑ��ɻD,�x��dlebՌ�7��ɮf�*>�r�{D�_��dþ�������j^D�^��{��tC�\
il�?�-?�>(��d��O00����H��̸~s�U�`�J��OX@ڃ��*�8�����o���aݮj������
z$ങ9C��2�`in�}���.��0D���Ҡ�6����%�Q��"a������ɳN������U|2T�9qp(�(
�b�V��h�mG��2P8��[ׂw���.&�`R����N�KN�d�7��{��`n�[b�T䑌faL*���א�����O*�b���H�i��P,��x���H���F6�Nq:�S�����L��x�	��K��0��B� B<A����%DO2Xo�Q&�y��S�Q{yHm�X4D��OL�M
ՍN�3����{^��i�)���D&z$�HK̂e0�$`]%m�Ӏ��0�VGn�4}=�>���~�(�mX��׀�@k[���z��"��)�"��$�}��oKIA�WH�ߔP���n��~�F��\!C���j�]M%)����D�isw�%UYuY���*�T�J%*���J�)���655�j����O]#��P:~��..2�!O�<Ym��k�f6Z��g���~�bo�l��5OaL���),�EO`+(��j�[ld>+-��9�5���f~�ynZ��"��\��������:2W?L���.5{bm�ǵ=�q�Y�D��ÇI��2Y��d�a�/{Cb���HC�����c��mv4R]͝����㇏��~,I]�N�*g4'T
)L�gW5��W��۹A$g��%`s6�Zڀ`8rw!��o>���!�5MZ��+���i�},]޽syW(��r���1b�h�f���wߒ�^YS�������4X��H-��6�T�c�Ͻ�s�ׅ���E��A��-j�=M[(�J��#�.|�Y+K�
;�L�U��8�O�7R^{3�e�������`eMZ�k�(1'�Z��/�H�%�W������^k���E�S0���iP;z���7|"�7��j�ܠ�2ElQ�=�^���2�����]3�"��%�8af�&�d�o�A�9�1���b�b��>�z�fd�;
��mծj�2:�[�y���3�~��˯H����&=���,ԋ�x%,�?�'�L�O$xn_���Z��H��|�rr���]ٰo{��>B�c��}B�c�J��x
���������j���w�o�<�*s>W\�M�BNl���d�h�9*�gD�����@
rP�1�89z4�&�bN�u^=o�[���j��ߖ��t�E��&���C!�#֜�\#_���f=������$�F�m%����)TT�΋#?�A([���9e�?�F��WQ�����ڦ��K��gP�<~|YpYiuA��u<1�g�P~��a�}C������ͯ�T����Dz��~�Z9� �$��Kk��BQ/Ǹ��L����u~�8L�b���'�@�u�R�v^��b/N�m���a�E((Zy�6a��r-4��`c�8�f����=�P��\1�Vȴ�O$S�W��3��o�r�AI{��hu3�K=����"1 �?�2iC���UI�;o�^�����zε=t�p�1���1��n�*2D�$��ГIq,�Dm�����)ޯ�4��#�0��S]Q�g[� ܛiZPei0��ߔX�Ql2�'�a�LM����¢���T�1m��P��ʩ@3^rVfU6T�Ev�a�Ј�x�.���e�<��w@�/��a�}v�y����� -�^��_�w%�z/�B���s�����Y�Tl��ߘ��m$�r����$���ޜ�n��+�\����_$yJE=���K��xM!���%}�e�)��\�H3*02�zfDW�'�0̷?t�>����9N[`�]ϯ&�ܚ�|�/�ͺX�jfrrq�[���O�'h��L8�C�s��6�%U{p�kD���P��a��|��	oR���[� ����1�q���+.�A�' �1Q���%Z}(���ʈ���^��P\T�cv}���W���z�Z4�� Dy��N%k�36�훘�����D��D��3%JJI_���rl�*�s�~j��)�Q2�����c:4Y�>[Z�}�Q��S쉡�X��vx���:/���p	h$~8\��������:�hA��C���>��Q����9��%_�����]�-3%@[�<Մ}��G�� �|�;k����}a�`���0l�1�wy�P;��7�v���/���v��0���U��Őוڜ25�����QW`��6�`t+=�8rn�6��5���a˺wa�Q��6��j��$�!!�jQ��5�����n�Dv���������K���_Ov��*"�����������#�L	��}R��T��eD�9��������4H�
�j]�5��8��m�Lw��>+����}��!�w�拗1�u��b�F���y���ұ�|����߯���	F}D��#t��aP���'������*��Z.��~!�st�ܵ�����Ę���ᓰ�f-}���A#��ߟꞂ.g�X��*73�hZ��ٙ����E���.���*:L���]���4�O[3�T��p0A��Pf��B����k��Tb?;�-��/j����B�ԅ�͝&�|����c���t���,w�9m?���X��%��@&�"#*C��_#!��ߜ��w^h]l9�o��g+�<�h�#��R(�_��ZFj6�da�*;���MV|!A���h�����9!ϴ�/�����6�A�? ��W`Vl��B��ɝiv���{(V�ˈ��p�#�-�sD��$3PU8�TP�Y��7�ȅ�E��:��Wף�-�Ho�nԮ2-�dM���:�QX���;����f���$����ްa��
Mϋ]��M������ʟ�5_F7R%W�T�Z�^���v�˃�I�3��/���F���:]=�Ѡ-����;���);�����Q�8�ZU�u��7���s;B�(��{Sj?����������𭻥��,��"��k�����2_{#����ݯ����.W<w߷���[�������k��Y4`�5�t����acT9C�S� v������{��B��E�z�ͤjJ�3%�-��߷��5��l��D$�a�Z<˿��۳�t�?�Z���>�M:����	��}b������:�3|#�q�u��� ���Y��r4��6���t*��ۢ�})��!� ������A��i��@͹��o?�8=��B�u9���9˴q��'�YDH��q�8J�R׭�e�ƀ��{[[eNL���?�F�A%�q������/�-�Z���nd�5�[w�����Ag*�8�� �����z-?��z�L�@k�; \�(��u�$ZH���D,z &�=�>����/�Ҭ�2R��)����J� �}I<F?>��k�	�O�kbk:9?þ�?���H��vf۶:y��+!����sP5�=%e&��v䛌�i!��h�^��]+Ƒ?���X�q�w>'/�6z����g%�� �[�@λG�uHA(���� �-7�:����(�Z����\zW��bRaQ���i�s=���ȎM�X �uY��*0�5�I�Sb��֚��Ųb^�>j����	��MZV	�=G3�CwHH�Q��rquS�Lq�!ɖchخs��s���J��/���G�>�L� �[�/>`��H�Ӳ}��ǥr� �3�y���9^�S��!��s�_��O>�ř2����������i��S݀X�׺�HCK��h׃�~
��ډ�����h�5����g���z��I)����$���Z��
B/�I g8�b��뗣���������S�(�� �q��c�غ�j&�q��@ǘ���댷���R�}`�֟=I�z!��u��v����hkj�z�u��
ɼL�r7&��l�*���3�����6w+�x��Z�*�&X�é���Ї&�w����f�R6oT}������/jj=�����G�%�@��1(�Ҁ�"C^
�f�'[��o�3S�J�t��3DP�#�x6�+�<?�TH:k��=��~���w0]���$�A���!�Jq:7�M�~2L��3�B堔���ekk��q�o;A�rE��N�!�a��VHo봱��TA�����H��N:|x�lpz���|F��-��WA�Ľ��_��9e��X5r�����"�Q�M��a���Y��(��_� ����s![_�s���?}��P�K��*ԜN>?볰׹�E�M����(GDG ���K~�X�9����6����9���Bg�M���8&/m�*"!I5��ͷA$��?�g����ЀK�|~!�ۿ`��e.�\�u�u��s���j��H��MH�����)���'��ʁ�<@f��:�b蔥8I��k^~e��(�>1_T�>@��������A<�2�d���]���	՝���s�J��Lr�ʥA�V25{����K������l�{7O¦�m�Z��%]5�Po�p�dυ#��Z��A��¡:��9m��$kز�Y�ܵ��0�9⋈L����1֢�^DGˠ�E�P���=NT�o.�d����a������ӌF�U��X<�� �3�O�+���((�!({`J+.���O����t]`�LM!�%�o� o`-�����@�T�(m�iMTB�˘ݢ?��2
�\��*0��`�����0"�z��j�����<��,e�r`4¾�&	A9B��q�v-����&Zx<��w���#_�*��e��ZJ::o���uQ�l��S��̼�c
��P��bɀbk/~�VW��J8'�B��D��5���kkQp�j~ҧ�4��AG��=ggv."�]��;t%Ua�K�a���X����_�.��Z\DX�p�
C8|���2��1+���}��W��.z֚o~�IBȕf���hk��*]]\iI՚�rڕ�$T䯀�BƢ���7s+�D�*s12Kx�	z�a��A�~J��q�a�$�A���hB
���a���I�_����/I���y���k���o����ށz���r�hJ��$������La��G���F��y��._�*�O~"�a���� ?�#ֺr?�P6t}��iӐ��0�rd��à�C��8��հ<`�%%��3��ȌʟXJ�Aqb@ sa��*Y������UQ	e"�C��j�\��Ca���Km9x%'���J2`G�'�aфJfQ͎�An���"�l�憈l��6�����UUU�Pq}&+��#?/�|/�Er�}�-#���ݏ�.{��'U
�Y����b�� 5b�����.�Dn�KK�\��03:���g���5�bŢ��K	��z����S��2�ڙv"���Z�髢t઩؏r,�lzY<�������c�2>�w��b��G/��M�%�n��4ds�-CIe���,���Y4�'2R#�-�)��U����ӄє�TF��)�%����(��|;�g�z������n�fz�w��Cmle�
���J(ن����I�����I��_x%��Hc���)�:>�O8ҳ���jC��"Ue�Ż8��ך"|6N��&z  ��L�J�O�X���Zʛ�Due+t�q�*���DK�8�RuSVP�[����;V��`���f$>��_��7��|��(ƀ�[�H���(�cŦ�xO%�8�����o?>
.�M8�XS��56�&].X�#��o��3υ�`Q��4�����z�L#�IB�l�0ܟ�L.ڍqT$�j�(��(ׄ?�*W�u_�{n���$��F�R�k���U��SC�e�4���33���6j�%���]�y�v�$E���!q�\�B��`i�O$7��#쾹��S��L�m���`���.M�9򈋘"��}#�u�+Y����~K�|�s0yc���O0�|��hk�3��ʺ�E��.�K 說������B���W`"Q�6f�pW��>�]oN^;�z�g�I;A�Sk���}.ģ5�P���i��1���3Q�v�������Y]�ӈ��9v�g�k+^�k̪�O�x�E&A��v��f\��������8t�O�h��X��&|]�[A-��v���y΢����
)�7�Q�oW�zh&����͇ƿ��~M�3����%���9��)0 �&s�AъC��O�]v 7n}�5�}ZE�4��y������Qu�+�y!n��2�8n�om�i���1���������tqk6
���ן���hh���?}�W��~�M*�;��v'��x�%|jS��Y�^����J��g�Ϯ�Ig��t�����t�����'y�J�2�r[�k�תGP[��~��H���iV�c��P�v����c�'[63��Vqܫ�����b�8�w���0Υ������)�j�n�K�2��^���3�������8w"��z��Ĩ��ϭ��@���L~�r~���+�����D��U�U�nh��!{]F\Z5�	�GWɾ��d�(�l�+���3�O?5�qko�L�wsUM3��,��
�2
ei��G���߼���J���*E���*��I��t����H�]�}����,�I3l|��W�P^w����Q��;�e7~����`[H�o������6C��:�u�8�X��䗺���vw$�E���լ��Y4�tj.�6�h�Zf��bv.���?�0z���S��;�ta���Z]��,�dq*�4��϶h�o
���gM8jCN:f�^�,ew�T�ss�}G!o�|ej�"\�rŰʴ꾑fzp�K�b5�����hnQw�Bz���SP�^Y�G7�J�n�ޒ+-��65�c�"�Ц����|�:��4uLK�cŚ�*b��-����O;^@��n[P����qN�%�����c��������^V�w�a�I,Rh<P-Ï�LMߺ%ȭوTq�~
����?�vz
�P�9$����e��l��%�9k*vX��.g�\Q�Cq������C8�R�3����,�{||�4߈���������f>���e*�^9�=qZ&����Y�B:#�����u����oK�l��̣ )�J]V6�����r�����o��.C;Ii)���0��*h�m9+t䮢l��8�{k*��͐��t�I��9��s��e)�u�{�UP�Kv+2Lл@(��e��gX,$�}�����B���H5��'Df�Ϡ�H3g�3*6��i���$��,jЃb3����1�YǮn8�6��<����=,p�Bfq0|2�!*�b3p�Ǻ�wqqqsKy��͌z�a�m���j$�<�C��L>�R	\Ԡ�Li�^rT����+9+6������E�I�����vJ�˵���%�Y���/Kq�J1��\7G�EQ}��*l���2���s���1b�$��A2���N�u7���iݬc�.N����5!PQf��Ī�s�]ϦV���hx�9W�����b���0�U�Pu��\%����Stȧ���C#.��t�l�t(�F�;�a�zYB &pk7)�����'Maԕ�o��W**���Ul�߭��_�b{�٥��.�G��f��L_��h���#!!q�ߛ�g�m��>)��; <G(��y�qg� ~g[33q�4}{���*������6�����G�lH�7i��r٤w��j!��!5�����z_��Qþ������*�xTY�Dr�IItb���C%JI3��Ŋ0(JO�4.z�Q���V�2m���RGSRHBb��~kk��o��d�g���#lD�Z�G;D��E���b{V�����e���Wa�`��N�����d&�����ww��M˼E����K�r�uk��͇�Pȴ��޷�;U
�g�gm��:Ls�1�捺��2M��/���^z�e@SW��no��iiي\FJJJ���s����=����X/|B0�ȣ�P��릝/-�v��Y�/��8������a���ǯ�5?H����3�'����9�QH���?���x)%e.uQ�Զ)yh��'$��������HEM}�!���0�ypp{���ͯ�j���W׿=����֊��x��G�YS�w�� �Ͽ�2�M��~��t�E�AV�?���C���T��4��������௪�߂6���/���i�*��}�4��k���f�NٟO��Y��+i�u'ώ$@@+fo���TQGG�������f�z��N^#�/$�ҲVǐ��2z%(؝�a�߼�;
 ��]9�J~	���N����hvK�Y^�[����U�vk���}�w����6?KK��'2X�<��O�r��摁7@%��(,��-^N��f�=��ǑQ��� ����+-�����K J�q�o��<���l����j6VV����;$�G��1Z4$���(@z��A��;�z�1�g#4_IT	��Qz
��Gr����=�R�d�H-�����SXGԃ+bi�쾬^�c%�_
���Vߡe�@�-�0�s��Y��3PL��f~�T�=�������L�F�"$�K�k�2#&|������z�*F�{����Λ^n:$���>1��$\�*G?Nͧ�
DX��plV����U�m�:�L�j�ʘ^JPO�02����������珫eK�+��Q+��6%�PݬfN�R�(���M�1(��L��N?=��(���FZ�g��&Ydd���c���w�(��{��G?��~y������
j�P7�����x+��jkYo�"�u�	�{���+��ý)Ν��"��:�ZWSKzD<T��w�6��>�_ű�����~�d)#m�PS��+%{���@3$�+���{f�yʼ��ڦ�m�O������%�Ô��WJ����y���Ȕ�n��kR��0:*W�:���8$p%�~:�m���X��4'WB ZYY�1zz՗��5�����{{]2�1Q�%1�9+O�|.�c3�j�s^6�B^��Ɖk�o�a&)��\��w��w�����^_�����.+�˻$�I�)fI⦽,ݮ��'J����<�k{�7P�	���#��^�����J�y���������װ������&8R�����/��7SVK�~��1u@��<��j��kL2G<Kg��H��i�H)ᴙ���,V��+uW����`�GP{��M�����Q52�G�M��mG�ڡ�7E�q�zӆ�-�����+u����ks�^�;�b��g�%9�*�����@U�F��)j~?���W4;���������4��]rR�N���,w��D�����S�ǋ�G��A[DulLg�SnT#�S�B��CW!�惷1��J�Õ3�*Ft�0!��E(��Zs)RRkt��Z%�"�=Ҙ��<g�"���L����wsC�ޠ��rQ!Y�4��
yXnH��k�D�+}��_98X�@��q譜d���MP��y����㩲#���<�K̬_?�6�$^��x�v�)�U@}{Q5�m�q���Z#%�O����荢���_Z��FZ���3
������ݻ��o{����0nR�`{� �cJ�8�hj��������YD��Q�=���d��˧/�n��n�z �ӀH��ﰨfpÿ�b/���:f&���^����[�|��b^[�F��԰�ѷ�5FD4|ע/q��9 @"s����������=v=3TD�|��^��]����@K���L���V�M&�a{�ɨ/��t�������_��R8������h����]���d��$�+l�R+t��;����:����C���'�H�P�|�ڥ���n)5��F���n��Q���\�i�c{���?\�[��Q턬ƈ7��8$��: 	�z��/��s��!�3;?�������c�2g�����f��꓾�F��\��<\(�~}U���/^��]尜��}�Y$�����<�f�����e\�{uC�����\ܟ�J�:��	1�����6c]�e�6������]Fr�^e��������C��H�������B[A6v�ң�9�ĕ�м?�{���QT��j<d�Of���28B�j)|�f�2`Ѵ�z8�EU_��.N�r
m���E�E;�<x�N-��tgz�nJ<x� ��&>fSUoL��f�>ɳ�g�?��ǃ/Ѹ��8{�J�z-����:��2/��y6y$�wnn0��>GR����/����x�{���Z��L���5}���{���v9 ���a�	�M��g���s]K�f��ff0G�a7@4#⇂���������G\)����/���PMHϥ�Phc�Q�C�*�u7���vY&>>~�s��m0�CʌV��^�h������>�m�E�.�� ��b�΅}�7�-�����u����A�
���.�'x��pq		�_�A'���7�e�m����޼5��g�Rb��TM��|�<�u���e�y������m�4´�^�~M�+�3�O7	�=�6E9�řޮl���{��^�f3��,Ͱ�!�c��	���L���l�}7Ɗ䛍��� �GvKz)e K5*u�|�tٲ�o�"��U� �RQ^�
מ��>}�_[~�A�3�Ǚ���q%���X.����$'����%�k�0�x=����a"�g~����u����Z�*�� 	ݜ<�ng{�ډ3f	 O�o����V���W�:9�n�)��-�͗��B}��/lƔ�� (���-�gd� �O AW�IAg�M6n�;2pssS?��Hn�˛Y�C+�Umڎ��f5K�P;I��������5m;P�H�]`�@@�~�o#���y���N�
�:l=9~�y�z�J����w�7���c{lL�V���6�l\)��2��K�L����+�Ԁ���v�:Z�~�����A��߄f�I��5�y��R��#�^� �������-އ��>��>[gEK���+��l�� ׷V��g�{�� �.��
�h�x
	I�'�2O^��Y�-i�^��V��6[et} hl��*�~YB��~&����M_��-%���������!�o��������>| Jo��yJ�H\_
���8�n�?�H�����
>����W�B$$Zm�5Ț/��ϊ�O��(�$�-ޓ��ʊ���.�py)hhngG������5<y�Gwu8Ylƪ����x;��RCC��ʺ�@�Ԭ���
��l
�V{ zY��5\���s��S����;��C�0�Z�6�+��-HHL\���M*�p{
0�����vY9��Ln����{��	�������<�7� �ѯCT��b��Nk �������rk���X/���O��Jm��u9i!nk����F����{u�%Fg,7��ɕi ^{�u@��A��@D��ﶼ�����ռ�C|mgo�'�ʳ��[&�kpE=�_�!�/z��������~�$`�����rVcef#4g�&�@�;-9�Pu������f�����Y�� aӐ�;�N�<�*��E���|�r��ޞ�_�"��s�7��m�'y�����7P�]���.��Dd��Lr�jŬ��z]�"�~�RQ�<�y��U}�����u�n��h2���?짪 �ъ��;\h{k�	���O�X��1�����fk>{���c��ܡ����TM)���U�f��vE����<d��?�g� ])ty.�KXE�ӈu�h抺�|{��m�zě�:ֱ��D�`*�#�U�3��[Z=3���o33@~><;!��m�7D�����i?xHq�P��y��_R�z?.�ߡ�v*��S0Zr����]c�F�G��C��>j��բH�0i�ڟ���v��Y.��.xо��s:��G��xB��_���V4!�X��^�a�����I�t��z��j�P�&�4i�	\i�Y�j�Q�aR�����t������ߖ��o]9N�V�pF^o�_���%+=��wۮq�1ypQ���ꊢJ�0���ߗv�k"9��9\���`W��	II��=��{N���^����wtt��U���	�0�#��g:����})������������p�f#�T��������Y}4&��pL�>
�3fc�u�������j]N�\�uf�����7���-�=��_V�����K���:^%7p5����3���ӘC]�.G��N��*6\��ʗ���]&�TW���Z�~��>���y����WG	">w���^�ƭ(�u�C:�~��R��}�$�[�I4���~��v�֢�bo���C zx�" ���lrs��ؗ��',x������6GPYmBI�����0�z����}�>�?$�����N��|z��r$9N$:�VO��b�C�ҋ���6R���C��ayY�q:T9T�`e0����q�7æ�L����ޚ�������r�}T�@�L�H�O5�	��N�q���ۇ��P�b������z�^d1����hiii��C��N%�9��q�~g[AG�肮2�7��=�@������,-�4w6dz�$�����m~���� {�8/��_�*q<�e||<)p���w�������H���+��Gw#�} �0hj��{u�A�3@l�`��-�T�s�E������-i�:�,��� �18���~��[S�a!@b6;�d/?�߶\��)n����+į[����I}���d{B� ����I��m}0���w�߷8�􄇇��H��~�x�4��_�I�"��
�ş
�]ww���ף���?\��V��>�3���n����
�1�So��p��#�5<�){O����BBB�,A���;?�7P���y@���j��� !��o�F^��oo���(�`R�4^�h|��Nt2��*��߿��=��<�:��F@Qpq�V��a%�,���_):ZbU�x*s|���������2��~$�� �Z����/�؟u����v�9�\N�o���<0ֽZ+��,`�a�!��y�q]An.%e3�;�Yݏ��o����ր��ylO<"�tsTS"X!�TV�iw�L$\�dj�[�7r K	�t���� `�InX���*���R��[K���\ÜH��{v<[TTd��gCZm���c�� ���h��昀��S3bב7���{�r�8 4��9���:�A����ڿ�o��Q�zx:��+=������z��O����Y `ќ�9�����E�]�ͺ|v~޶��ܲU���ƅg�+1��,�;�L�Bf&T6o^��!6���Vql���6���rBeŮ<�Te�5��:[���p���w/s�'����r������ׂx����ʛ�>�����v��w����]�#�A�'�����?����jk���ʤx ��#2��5�Ԁ!y#eee��� b\Do�dfe-&���eFI�3��/�}��Q��+����?~qq�l2..
�٣l�G�H��W�W��ueI!dgG�%���=��^�޾��?�p�s�_����x�s�m�'��+
	�F+cL������=^6t)��?�0���S��}��y�v�W�qir�
����NT�*?����ښ}���9䐺0V%G3�C45˟������))᫙�;\}���\[����45�p�/�/����1$��z���L/�V>yYe��7P��� �� ,�e����O�6�Q`J�K�S�G��)~4��/;V�SR�}�w���O�~��Dt,��(�SSSn7���ի��ΟJ��n������`qqq|�V��Pֳ"	�M�G�{o��Q{����<|�X��w����b�P�5�b�����'�i�������4����2�(�/�sLtu�&�X��a6����t�]@ծ(����+exݝ)�ü|˳~¡zj��`eu��*bbb"U̩�����w�ƉI!���<�
f��������ˠ�On��r=��.2�����_����U��2}�a|���h��e!��TQ�N�:::���JKK�+�������4Iuuu]���������1m������rH�c\���o�7����w~�5�&//����)_2�����j��	qp����QK�S�$����[�U�`���}������0�'���WP��"��5^�� �]�"D݃���g�	�)d�al_��-�O�����I-o���������$�J�s�t]]]ww7`ǉ�J|�lI�9�s��l7�8��EE�O��
��Y_e㧉�07w��u���?<___���~��0}��/�����5a1�ŀ![��_��4=��yWW�|����վ�Q���]]�h����>��@j�~��?�Ƭ��\E�J446�W����^ǇʛyxTMm�qs��*�E���<�2�@��3�h���dm��%���ͤC2��`aa��"�|�{��5񣦱53C���Z��kr���9����{�.)	�q�7�c�&g��Rk�<8m��<�k'�=�W��-���77�M2��	ȴ8�\Q�N�zz
KJJ���"5���ᐭ�	Ĵ��F�:��t��m\�+L����G��p��7�oE���7�]~�=)А[<�"�c�k�c�����5�q742�6�(��S����`���56
���w�b��ꎵ����|��*`�������i�y&2�wh�l^���? ���!' �������G?b�ge573�*/w��l3X;���T�D�4���x�)7aQ��Z7m+LOp��\\\:��&a�����ٳap���"H%����ф��j�p*��*�./^�pt,�ە	��}��2��L���d�œ�/_�ς8һ���Ե�+�[W -�y=��Z�L�20` � ��̀�ģs,_:�f������q�/`�0��Ǐ�}��-;�#$f¾����
��Cr�VK�T��%�R�վJ Mbxh���f��zss��T����gu�i-�c X@ׁB=e��.�LP����LEYXX���/8�'ܿ��8��͍?l��������-������0]$.8��B8OP�8�ĕ������à��Y|�@]�����g��:;;�k���jW����q�#��@�"��Ծ�`���::�%���nokO�7�q<>=���P���e��<Lȸ�"��k�NQ����'N��Y�9�����0��}����##:��)����{�ne3[YY�v��GR�����=��y�+�,�%�Q�����8�V�����/��ϹH��o���---�(4��?00��gFKC��g}xtt��7Y�kTfB6DKO�F��"����f�����X��8��1@	9<<TPP 'uss���((( �x*۵@_J���j=�`��#��m@�%߾}JO���������D����`���ɴ�JǈB[?~�(d�/,,���8��}o^�\�w�ם���c�u��� �]��5����.��b����e�kYh`���w�������h곶L�K�;E�3������[T}��Y��d.x>O�E�[c3��.(,�~su���822��O226vzrBBJ
�L��ݻ�::9����>|��<����%;\�4�E�Cٱ����R`��K�।��uws���DG{�J��\��+'���AX?C"�*d�O<��&�.$$�`����w��"�9+_�[��A�rjj�Uj/zYs�@xpw�b��[M�M�|��,9
�[[[k�_�ǿ::lll0ړ�))ty�t0h��a?�F�v)�&��cB[��q����j��^�zO�o۞��5So}|�k�v�v/�M���*��������>1���u�'=�n 3���[��ɪB��j�)))���߁b;�tV �C��媓�bnT����w}����Ak(@�g��@���p^���)'�d�k2ͣ�Ʀݟ"����y�����h���Vn��|0�n�����﹙�II�,Ma11$�����AP��� ҜK��2��DZ���ʩm��4;{{�hEV�w���K��ˮu��� ���9�I���E"c����=2�́�⤲wtt��K��Ѵ\���4�;�Ô^0�@%��-�_poaW�8P(�������+&���}�_�(��V��p8�l��Wg�t���y��lD��>f
�rIR;a
$.;�O�L�jB}���uw�ӧo~Ά��B�Q#L����+�p�A���D�万r���כ��ujkk0��4eg/��[�	,K�d���m� �9�ݣxg�"}OOO{{;�~��}�N����١"�LS %n��,���LM&��!ƨ��:,�.y|2��臘�J�VUU���MA�g�x��L���<�?f��<d+�/�:�ŀ>2��_���0=�76.��<��i\p�ŁI�ⵕ'����a9ͼBM�fivn{�FE�n�%������!�ب�%�����.@]�KM��L�7�w2��g\o�@�}S��W���7/'G��+�b��t�d#@F@!l(o�,�K�7=�k;t��0�t?��@���
�7��OSE�zE�ļ��3�S�W�!���9�@z��f���]��5�0o�`lSHP8p���(��A�67g�A�X�W�l�QHX�M�w�'s{artt�g8}WW@��94H��2Y���f�̏[���1������9[������ۛ"BL�F��r�0؍�͎_�LYxh�SR
�㉉�Ef�#rP!��Z�<���'-�����7�b�||~ �,+���W}Pҹ�k�?��_4��s�@�ꉯ^�V�0�F4Ƅ�i��Y�=�(m6S�#~�څ"*۟v�<�,�'��
o��~$s�@z���߿����CRR҇4���w�&'&�ŝMW��/��	�M}��!���sxp0b|t䮠�����b"L-�����lw�{�ή̕\�,J+�����")��Nn�Fg�=H�Z\Z�*T� )�Z����8s���y���T,G�@�{��SiS���~�"k�2N,n���%%P:Z��o�n?�>�(��T���������@��ƀ��ξ--*��K�u����������*����6�р�D���3�ro��/c���� ����t� P�6�*�\�:��������vs;;;��vv�����Q��ZW�qu��L����qZ�w��ruu�����!)!G��1�s���E/��n~~}6~��L�.Pa8�ݭBQ�9؜�@�@��L������$%%���NRõC+��wY6�i��@>�/`���>0V����%ӑ�c���|��o<���8:D�션E����pLă[������Ʊ�5S��uCcc���:�KN{��]==ܜ��v	�<��	���]��%$R0[���Ĉ�g�]"Q�� 7�L� �x�I��[f��[�=C}m���$=a��[f������-��-5��vS�GL����(�̱M�i��T��	qq��Q����_�G1A/�_�Z	�M��3g_5�ã���Mhh��X馻��Mc���;~;�l�r$����}���;�����!!&���\tO��f�4�$c��Y�&A�$J��s��+�G�������|h1�m_�+=��LLJ����y��=�E�VF�D!��Z�		�W�Ө��F��àA�s�ī�OHp�{I��(�pp�%�Pd���#/|�°������w` �ϛ7)}�nu�?�����񉊈���ccþ
=ӵ��=Ln��ڝ��_��VX-w�ϟ?�Har(9����F��<����uqՙ3��� ��9�)�A������^�(e6�8	L1�mxx�����I��h�:��(���M��Z�ziqq����jѦ����3燿��VV�ih���A�YY��-��H�$''L!n5�iL
�3	l"�}���|o4������/���R8�Ij�]��z2��6n�w�<E"����k� �����KNh��D���7K�#�|HNV0�|?�'+�]�Z��������nlDDDT���4j�����o%%;@����h��Ԃ.��򬿽h��ܩ痖����-�����ct.���/_�秔�W����j1 -�A�!A[��.��Jgi֚a�@�S�<�7F��vd㔮��Z..6
��ٓ�-5��I�[XZzzyc�W�H��� �@�y�k;������utw��Z[���03G<Y__����KC�8ט�b���*�0(lz\g*��8H��ǌ�<ͫ���E�Ծ��^���U߃�D|�Q�3��X>��ui�(�o@�\\\��+;��0.���W*��tn_,!S2ed+.I��l�@p���"H�# ɣ1���{��ӆ�-���E��iU#��׏@!4���vOe���cen�����5 ���KG�� ��z�VZ���v�q��){y �����t��T�@�Wh�a�����#1��f��?G���;ǃ���ŋ��<����4I� \~W�╟��JO��\���A������Wc%3un����r@^�� wͫ��:�����MHH ��n�����ZwW0�Y�ç	]P�,�6/�)����k�<���xno���<{��P�,P�� _k��f�1p�J���>�S��Y:8�6-[������ϲMP���u�x+s|�fea�j$�Z�Ry\&⋅$�l ~�wc�l'�� ��uv���DF�d��+����mzzѧ���w�H
b��F�����Ɗ���.�dR�n.��L�z/(L���r���ITL���Z�r6�\��۝�:]�7�]�7 �f꽜�F�A5jg/��K��g|�ȉ�,�ݏF
�u�0�]�MVgO������ax��ل>�Wcc�/_�L>0=B0����La�)B�s^~���J��+Sv{��VX�����<[T����,�Mt-� �l1��"�K$9�󭗙�������ɓ'��Re�mh�:��XW ��q�HO�)3��d%;�ZUS��e{����W�� �۔�NHph���{����6�r��j�ƥc�hy��`E�VǐF����iz���~Jr����oW��SԹ���	L7g�~9�@��/���e�:S������'��X�7��d�u2($o,��012�4�9�!}�H����������3B�y, B*ҏ�Ł��o_V}��g������F�inn|�$���Wn�A__�wo/�c ��""������c��aod��}��<>UU�<�/~�C�!�a ���V�����s77��'�Ia>B��y-ڃ23�h"q��DS��+�뵮������ ��3�[#ܻ��~�Y��d�6�� .�e���&�k�eo߽���e/�-�Fe����TʆH��0ᨐ�#u9���g���̃Pftj����aQ��XM�n��3��V�>c��S{q����/[g|�^�Bp'����r�m~8�� �5~Hvf��ψHQ�c�w���Oѵ�A���f?q�m(��cw�8��O��:�&A�]]��X�ٽ�Y��Ύ���0~R�{���p,�9�OR�m�w��g&S?///+��&~��.˘��;���棦��d��/��4����<ۺf��Y�X�Y��odC�㗸��5���o��J��O����� ]������|k���z�cN�q��%3�������!V�����B�X�c9���an��> �l:�v�_�x���4tRI�o-��V�����orw�_�4NN?������S%�J����
��HVz�+'�d+<	��[y�,��eIy���������^�Um�B�����fnn.)%ef "{B
��ϟId�CCq�{rG���Ӹ�-Z�޽&�ONz{C�c Cfnvvvt�c�3�J�!��+�O�03W��7�[[Ej��q� ��ܮ:�{>@u4q�g����Õ�\4yo� p}__��GL|�R��y��zVv�j,[����՛�&�\����L��� k��Kc�!�b��p~��Vuo����hj�A����F��\�N,N��X����2�ӆ����-�W��3:;a���9yy��>A�+��������lʫ����ʿ�i� D��3�L�	��=š��h�<;2�cd43Qa\�߿Q��h��3/�+O�-,�Ɛ�0��_�qq�	�Lg<� ���	���y��^���ٟo�&'���'�����e.��"۵55�z�u��.w�� ��ERԡr��� ��=����@�oؓwqyH��@�٠���K'�u�'e���aKފ��=����&''/./��<����514��s����>��]H�����L���f^&��8L>�����
BPPR��/�8pvv�yw��t����&e ƻz�q�6o>�H��Q;��(��~�Vl�y+��22�{�)�A|��|k6N?A�E��J��$J�a����^
{ۊ��!T�f�個����XV�ɕ��UK8IWf�G���DN��}���tfiN��@�X �j�<4���J�n|^�.�zua4&}��.ٌ�e]|!�Z\�H'%��l�>PP а������f��50,K�	��G���|c���?�L�J%��
���=< $�Θ����/�<��***���wAcPK���H��='>�:��<��g�,			QQO`|��HC3}����x�J�~�(����53���n>|H\XP�7usJ��Ϟ`�������[RyX��������A��}�w�z<FFF-�\\�>'�����G/��8�Q|��_������OKA�i;FA�E��o.�+�[1�ZJ�	CsV�z2)	�D9���!j*���d��x�2��a�%S?�e֔������I0A������4�Z'1<L6�k�!p��ADa�b� ��Q�#�ej�J$�;���,�؈�E]5�`Q3UXX8�.u
��.���1��r�B���A�p�2���o6��x>f[;��81{ �8W�v��[V}������ƛy�(��#[_:F$��&�6��
�XE��+�h �c�g�1quˆ`�:ns/%*�Z��a}vj���|Gs�%	��jw�/3���|됯�Cu�W𣚱����>kv�����=q8$��Y���0^�f+a��!!�a��`�!vz��[��@UО��c2vX�`CP�Ɣ%-g9v�������d��5����\�_�w]�����}i�-v�� ��bcc���R9�� ���C�s��?�����)��9?MB멪�]�DDD*zxS�"?�@"9�PQ�03MR�����𪊛�z��N�}��r(dZ@}&8v�}a�{!(uPe�c7�3�s)��'�C!��R[�G��K][��A��N��2P�1䢾-F��h����/�B��y�j	شj��l��zf��~	�6}�����V�u�Q��/Y���h�����V��-�K9��>�����-�2�Z�j��$� �i�Yԧ
�x������!1�$L.%~�}�>�NcX&Li�V�ٹs���1��ip&Y�ն;�3tKU	�X"o�PK   ǕeT&č  ��  /   images/dc330bba-b31f-438e-bca0-f858f4ffe113.jpg�	<�m�7~���E�mDEɾ��$I"�RLB�$[�6�d�B)F�V1R��/�Ⱦ�1CY"3af{O��յ<����}?��}?����ǜ�q���w,���{�c�#�I`ˡ� � &^�y��9 ��v �� � X�	�y  N��ay^�k�?��;��oǁ��?��Y �?����Q�d��?�@�ֿ�9�� x�|_  ����m3m�ʹ�6�f�L��&G�����dm����e�ݽ��e��T�T�����U�u4����Zjj�jڲ�zZ:�Z �}�` +xR��7�"Px��g�:�:(����8TM 23/�v��;c*d��UBgU���_6,�d=�i3m�ʹ�6����/LE�@C��;�+�`��;����A$�e!���a�؞�m�EP��已�W�3{�����8`p�����8`0''�/77���V~!i	�������vY�=�RR������kii���4�T4�46n����������&�M�_N�F@�lY/�`�@ �V ���#��y Icec�qprq�j��C�,�P66V�XH��c`ܦ��}�QW�\��FL�]�}O�����k�����رSAq�n-m]=}���,Z:f����I'7w�s�^�>A�!�.�^	��-!1)93��ܛ����/.)-+𴪺�Y��u�-�m��]�����GF�����O�gf��IߖWV��)k�v��[��v	�v���BYavAX.oT`eۦ�.��(�5`��F�о��O�8�5��g�s�l��� m��òΰ�˲���n��'� T @ ���{�\�@�gk�n�R۫�WzD�U� z3A\@+�o���Eg� �5���?�Z���F�SNK�ҡ�H�wQ& u!�e2��	D���/�2��d뀳�a�3��"�(�vf�ha�2{J7~t��I�4H��b"%ES��fĬc��&�fa�q��@���E5O�bg�� �9��	0���m_���Iv?]p�}ꎥ�>���ޔM8���1���n|�e.KL�-�`�8$늫o�_f'�-o�����0����E{��ESIbJ���~Ǳy'@��s;�g�T`\U�{�k�'�/�
�����w��%է���׉f�$�d2���Є�/Ҏ���>����S����G����ѓ6�y�پ�����S�w�����=�q6W��Ԟ�$�I1��E��|"�y%v��٢��X�����6R[,�w�؍�Sg��<���Nø-E�)��e�j��&�}�O��x-��
F!���0��s��9�~�^S�۲co�I�r��B:+�/TL�y��L�Wc�ד&�rم&HZ쳶{+�m*�� ���Q0�-W^�����+�K��ċ�}♋���g��J���܇4�}�Ţ��;����ی���^��G5��M�7�ϔ���U��Ɋ����տ�^7���ֿ�~�(��[��[�im�z����6���/{C�u|��x�ߏVa9��S�9*7�.f45wת�ҷ�@��s��S�s�O:�$�ڒ�
�$�-T�ĥ|�O�S�w�&rW�B�����>4�1=*�i������~��w�$S��߉e=��J~=-"�WZZD������E��mڲ^�ی�ǡQ����C�4��L�����ϡ}NE�����1
����b�
�V�ܾ��F>:O�������/�i��\���ܝ����+T�Ƞ��Bʢ��S��U�2}�	�`����\���˓�]����B���e8YA��pL`_!���Y�(<e�T��y��~׭�i��h!��N�XP$�q����G����c�*�5��+�w�b��[�QL ���:�.�'M��+���.��яx A���+B��?���'�:�x2�nhg��"��n���IC�����!��C;��>���793kl���).�62'Mv>o�&�܂ZG=��p��y@4�p�X�N�`t7:UƘd<�~�{��?��*O�k��w/��<�{A|��J,c��ӻ�aq�Z��Ђ�Aes�y�o[,v����y��c���u`��;��E�V6F��裦R��9�X]��u/��{W��[-U����:�!�&��!��i�ͧS���!H���5����q�1��3����{�_��7�5a�| 8���q���S��'����i��˰u_��b)Ƚ��c*��u��C���=i߳�2CB�[E�35��]b~����q=̢Ә�ĩ-Qv{Y�X���!��#l��s"��:N�g�d�5N/���A��8CvV�?��۝fr�!əe\�'8�iP�������I�/k
8Y��6�Y���.��.�J����m�"uf����ˆZ�3d�*�K��픪 ��ڒ����E`�E���h=����O��`[}�ر�R���T�(�b 6�-�tm�~���yR|,�����u�kNT+�S��I��,�?pѸ����\�v�e))�Eg� ��)��%Sҽ�<�e�"�T�b� �e��}j���g3�����"5����	�,�վ|֠nt!�Qd��<��k3S����t%n�A��~�:5�q6Z/�vX�(�	�:�e�Yщ]/��I{�}.eu���.<��}�Ѝ��K,�s�`��6 D�u��~��՞�����q�e�l!�c��]B��mʉ���'����K<>T�bVE��#ˣ6@�����j���]��:X�=.j_6���yd���N��s�9/1���hb>	1��}�p�T��c-	Y�n�ZG�[6�k v��B�?[=I��7�:�=c���R�g�7��Q�e�V�=��34
hq��*��r���VO�_j:��xQ� ��բ��>���6�m�ݶ��9�`)��hMx�wA+)�pV|��|����+��ٝ���ѯ�b����h=�?͌�u���>�����h��_/m��ݖ�&l���h幰�C�����۟����6���a�s9�Xx�����e�jPke��;�/]�Y�B/]�Z���6�V�W�b����^����9t������ьF���
�����rB�OP�1�w�3�e�J�كL�o�Cx
+��6,f�/���=d旟AEȖ��$1?&��zd��YE��O_�[)%�B��y�y�⍗/��C������(�~�����f�������%��)�5�d�G���<�P� ��?p"��j�!=�/7����L���X���~!�7ߏZ�|jnzq���t~j�!K��눃0��͎i��Z\�ǎ�B�ݿ6��K&�arw^�BYry�H���rN=�u�Z].���h�;�˂Xᜩd������dέF_O|uq�,z�WjzǴCCm%p����S[�{�Y�����:��<Q�m�un��{N*�?��IوS_�K�C���ɧ�.���S��1Bv�����.���6)������ i?`�Y�JRMB�%b˫���X�~ڳu��<�-�-G
��/d���o�.�-�9)��U^(]|�Y�h�f� �66���q�yZ�jK�p���!�`�΃�!�zm�>a�i��;2�l�c�zb�1��1:�|޹c���n��9�����k��W��\�&�s��Mg�d���{1ͷi�S<<�:�{���V����O�pSG�,����B�ꤥ��v���·zN9��ߙ[��o�������g�XjW�"��G���(g/�ֿF�v�5X�����A`�P�ժ�ۇ�kJrH]�[-�#g��v~ĩO�i���ŷi(���h��µϲ�}��3��0�Y��>��(WL�|�=B9�$8�-�=�*;D6c�_�_��3<��fuHz8�o*s���_l<@�@ƭ�"nbJ-��r�~�:s�N��n�nu= ���}8����Aj-9|ʯ'��dW�ZUZ��߮�+�A���Q���fj�L�tev�Z�T���D���8��:����Z�7u�� _tV�L��?�T�X(�p�<x��y�}mf���l�s]Ml���=@���߳�A�//��3��n����.[5���n�󩔓�| ֚z�M6��tig����_Q��i݁icfܺ_�߱[B�?��]F	�<�r���.m�_n�S�N�>L\�s�T�ږ�Yk�s�)9���{���B��^n�q���f���x�+�#
f��8���?���8�7�WKy�%���ȇ}D����ഒ6�ӫG���zdMmJl�YN�l{�k��K4�@m[��^is+S�7�o�Tw�ɜ�kQ�Ɋ�%�lx�G6�s�u�xL�[�l�z��%�f����A���,���J�CJ's>[��n���s�i_��{a��+���������y���c�&β�n��:�3Z���`���}��g��l���oE<���k٢t��T�MG<��Z����u�
B��'�'�!��rSu�Xטd!"�/Zm�j<<_���5�1�݇u2�oq�c`5�A��u��Gˣ]�"����1P��g��"_+��NwG�:�{�^n}�g~�ڇ�VH�;ѵ��5����^P�.}��4{������M.X�������B�c�a���C��^a��_���x$������k=o|{� /'�u��������ؽ�*.DDHԒX�1[b}Nޅ[;�o2ۮZ��]l{� 3�Z6��$S{� �j_]_���ޜ\(�m:��&�*�}�-y���{e�T,�֒���n�_��5��N�c���}���4����yw�<�aoxh��y(����7�m�O__�sI�-,pF�WI}��s�-OS��2��c�"��~�L �E]Q�d(7�6�(I<{��T�>Eq�:F��:V�Sq��Am�Wt�I#0�eX+�@y�XIo��~�	s����E�@�Xm����:W?q�L�h�o��F(�-����WaL��1'��%�ғR�iK�R��Q�g���jE�_m�bl��;|��uyj0��2,��M����BFU�l]P��3D�m�W��V��_��I�]/���E:��Y�,�"��_�4k�Ʋפ���3��޵�%��X��m�Uh�l�����9���ߠ���=�V$;�l`��m/�����M�?\>I���x:ϫQ�߲&�ܸ�Vt0��[������Gfw�j�a������������u-���k�+�G�0�.8;�a�V���c�S*�_Ǌr�=�ŏ�� /�_��}�B���w��8g��gh��!�h��p°!��*���m�ᘋ�M�A�u8�����p���Ȱ�@ޗf�>i��I�V/�5g-���'�� ���;�����\:˙0.L�\r���F���R[�X��"KM$@=�8�>hΡ�qj�-�w��V�M�3�%Z�П�q���믋��fQ�)yą�4P��Xw�\9���p#k��^�Q�F�#����k�I�%`�~�C�2�]�o�n��p�;xs��=Z	�;�]�R��n��4Z���շZ�=BMʸ�����B>�?r��7��ۣY�,�_��\��O���p�����M5,�:��L)&S��:����a�{%�7����|�bc�RL���q��OF51�	�=�P�"��[V��nO��'�=^vr�4C�UxX]���z�k�7�;eD'4��a��T���Vv���WQ�nL�Q(˰�l4K�+�ê$�|�#���Sk�`���C���/Me��u����}Q�v��٥''���{~i;�����=h���39������ǫ<x��4�R����n˱C�{X	5���9&0�x����h-ʓ}�Rˮ�
�f'�H�|�I�\�ШyICu�� �I��i���YP�-*E��.����?��46�T2��3��������y@kV��@��_af���l�;��cw����Q���g��kv�;1���	;=��|��+�W
yZ�tӏ�C�x�����];���?KjQ��cA�U�<ξ�oq�5u��}����G��ܔ��
�_O&��.�JK*�y�N���.��cć垀<�}���88�̟>{v��hn5�Oc��trM��2�,r&��!؏��y~�d��,}�u�p�6FK��G���÷�����w�=n:���	hְ~Oİ��:C���k|s�կL`]���m5Υ��Q������l�����Վw�ɔD뇐�f�$���;~׉�(^XuyW�{����AY_UC���j��ۯ3>$nO}|�l�J����9}o�Dv�Wf��j�ڛ�>>�rFOE,�����z��~�������?�w|O�p��qة�|�o|�ɫ���ӃG冸��< %�TY�,�u��t+B�[tK֭N�}z��|�;޲�SV�� +�ڢ����.�k��������v�?�߅��H���\N�r��S	yӺgK!��yݳ �"�a�W�v� m2�@\e�{*{���Ov*tP�a��,X��IgqޑVZ\R�X��Ĉ�d�y�)��
��ɛ�y6[!u��/4�`�ƌ0H��!`�rE�?�a��9����U��m3u�.3L<cB$��O컒������e9�ـ�<�0�?eKt�Y��h���ʒ��+��W��ś�} 3���@>�4l|��l�Q.��;'A>XQ��K��!_��"�^X�\��K+*q��"��ht�+e5����=��{���j�Cq	��Zp*.{�'�~%p\�R���79��!>���N9w&�i .��A�e�&_��'���*�܏��<h;`��P�D+���zښ5�!϶� ���;�&�\���w��3��9���5�4���(�|�s�8yBd=b�3v�����_|{*{��)���-r��G.��f�����=�p��U5ħ�R�|�z/[���&=/�k���V��`���q�c�9=�7��/�\O�d�>�����E�n��Mh��|�`WHũ^��cח��~�o蓃ы�도xb��*�l����1�����O��o7�c�6}�p�?��~�X�u߅`��g�w�>�s;�U�bd�vC��w]x�.AI����  �ӐFƞ�%CK��/��M���KtR~��̐��>T��߇��<�|����}�q����:seN��|Y�l>�Sl-T2@3~������}Q�������Ζt��t.���O_��B�|��3��ӄ�ላǾ.��m���W����=0J�� ���o۝浣9����n3|���tv�O���[x��d'������M_Yri�뎴5}7�r���n��d���6�z�#��U�b�7U��e�Ox~�A3�3B�A���,�I����/�v~64'�Q��Ko�seH!k�t��؊ F��.�k���-�[��!�R�L~]��3�$�,,�	D`(������4+9��$�;U��s���ϡ��������� �>�|�@U�B�����Y7?�P׋��*j��"�����G��YO��
K/�
����
���j��<���z;b���ﮀ0��2
5�����*�w�B�A��܏���êr&F���������X�׶\�|Y岦��������������2XC9�ʅ`�P�A��`�G�[���`o���]���˅�x��s=�}��][�������������������������9��r�5���O��� X��,��5�?������?��G#տ^��}<���d��j��j���}�������_����`�go�]/� m�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l�l��������q��X����wBYX6~��
��ql|������������'���O���{����B���<��b"Bb�B�B?�C
^������)���+�/��!bAA!r��!��������d�l.��%���@;,�K�$,��p��+�~���x6�>��e"%Q#�cL��9�X�z��[K؅�!�[��FC����#�ȗ�Z�����qS	41�	X�")�L�㞋h�)u��ew��!VI��^�	��&b��CB�l&��N�_o�┏�S���wTi�>!�T�<8�*���>V���'��0v�|������h��C��I�Y���GvG���Cgwò���v&p7k���֊^��ф���|h�ؼ��邨ޮ��;8A��O6��F�x�ΌT篧�����&�{(�p�{��$q��XZ1�x��3��^���`{��"T����`��d���������5�����l��*��������լ�[fĻ��j�B�^~�N�u�\	�v@ی^\1����4����%yM��Y�vN�����~�lBG��Y&��aX��b �L`�
y]�2��82f�	���YF�1�3�6L�<�v��OKd�0��@��Qs@��d�lB�<CpQ���!�8H�IonA�5�����7l����5�ڦ�t<N�\���7���Ʈ'��T�}P�;�i�>��h�����}9��{�]>d����	[����}B��������6�u����ۼ�rT�I�	L��Я��.c*N�);q��W���t;F�j�{����`3�ޛ?By2���g��s[�n_CL��w{�ʠ�>��%Q=&�Y-u�����_~"UއMk��/�b-F��h3�3���H7�|&��e�����#�aʱG�ת�v�������L���(�P(c?�5���W@tl���hVJ��݉_﷼!����aWv�����&1mN���yA�7�����{U���Q�Q-�q&���E�f��L�S�>���޽4��C��2B������2輄ҧ�?�\�TFWt�C�&w�5����K���9J�5]��ȧ�3q�W��#a��$����_
f?s���j5�IϾ���鶨E٨������m!L �텄7H�PZ��#�ƛ/ܿ���$m3���]ac�.גP�u�E������I�~B78��֔���&��*�[���|�L�p�V���	�8Ľ�'Szaø�E�I�hiK	�]w�~߿��-�3��I�`�(nL�m�2I�]D�@-@���Ō��9w��O��㏐X��B&�>˞_ʗ�kh�J7M�i&��d����d@�3տ|�]P�*E���Iu�NAMbY�����)^O�+h��5�N�-�_�]T�Z7	�h��d]�G�L(lD&��Ç)��\�/&(�����c�ֹ,=�˸�
t=�'�x�:&T���)p{&�J�
n��(�&"�00������ 8��laM}�&�9J?a&F�GQii1��v��z���;��kc�b��]<8uW|�wIّ�C�蹸�ڨ���X�~6���a*�n�Y�ib�� ;&�������?�}x^�UuM~��I�(g�o�-Z��-�ꏓ�̮��f��y�� ��."��v�*�{�c��
'`�H	�X;Q���xRqyp� C�^�Y[U��'#�\Sq�=�T�{�ߤ;&��״Su�o�:[�>�R,C`�j����w5b7��(�h��k�q/��z��H��P/��W/�P�Z=)�'���-�N%;�H!B����+�3�!�0��6�~Gቹ��8��A�L�GƲ�40 �"��������r��\�?�j�Ӛ	`p��X��SP����c�~��@�vx<f}FJ��0[W3�/DQ�ZQ��ֺTM�1q�8c����n�LMj̑e䓎�1�F&�B��t~����o�%O�)��o�e�^+T������d�)�SGZ(��ڛS�E֦����w"�K���	I�G���%r�W���}�6p�`t!IS$]Fǆ_��|�� �˭hq#a<j�j&­p�`G�^g]��}R��o/��R�c���k#t��É����t�I�g�}�ϒa2�?7$�5 ��l�+C����&���D"�ib���PBm��죎�	�>�a�)Ɲ�#�ڼE��
ˏ���ޣ�LDp��6�vo��4�5�F��o� �]-�؁#ZG:�_'q��k��[�@�X�E��Ӹu�`(�|��ڦ���"�j]p�l0��Zv�3���bш��܎d~ojP�7��ӳ�~+���j�x�ہ���$�i��Q^"���sl�J����Ҡ��T1
��A�X�VT:�-=6�ǉ�4��E�Q�`TP:� AOEy�B�7�B&�E�1���ڼ����MɆz��eЕt<zQ�8N�Y�. ���,�]���3���=�Y�G<^j��"��_7�Z:1Ww���X]�PS��:�����]\��j�z9%�����=G
�.@���'d�YS�y'���sa���e_�8���E�SWz�������f?$#�O9���G�Դ� 
0LB]�u�'����VY���ǵ�)]�r�=_� ����gij2�%����Eӫ����y?�����"�>�_!��q�H!�9���GG�~�Y�v�i��o����!8m�$��(���;�z���)�k�3q_�Uo@����,ƾ����mF�����Fh�<v� ��W���C�
�W��J���q����P'��?�+����a��cx��mb�d��8(-��ST�H������h>7�1bz3��G�/U)��̬9(�5j��P�F���\)�Z9{�J>�7c��b4�䒎1����dm�,I�4Ck�=���CSxn��0c'a��r�cl&nOBb�4��Z5�}U��k3�+�g& =����t�����p{��=�e@L9�cg�-;�	H��T� x7�j�2J)�bS�q�f��h��f�$<���Y����a��8���W�T��`�[g�Gr�5����eZ<bVɩ8�����z��*,�$qD�'Ь�|�Z�u��},�J�RL��ju�B��X�q�~�D,¬�f~�@����E��<[g�*�"��
ʈ�W���à�[�|�|���	�'�*>p^�
������>��t��O�A�$��4z��j��2�����x������I��v5b{(����V�������P�#�����/�g����@���}��)6�H)���y7� @��z4��J�(se[Q���ʎ���d�]TP�u�i��e!��qP �u�&�<�'T5
��^�� 2�GG��C���+}�>A���J�����/�I�	6�\k�cJ��@ej�|�aG�נI�g�=��D$���T�5�sI��W�n��Q�֞d�� �d!�s>�f�9�h�d�;3T�F�e����B%I8&����6'�',��h�����N^N���s�j�_f���J�����2�ƒ�B�4��yU�#��G�=eF����J[Iܓ��YQ�ܤi"U�_<AJ�S&��I�����E˄>겛r�12���vήu�A&���?7jc3x ]>o�0B�[���=#�2C¨Q�A�;(�$�V�9/!��^�>#�b�l����l��ʼ��tr�dg��S��O�TUF�:l�:�lӎ&��q�#��=�ya^z����{���^�o|��?�O�&Gl+mi	KO9�c`�աֹ�ĕK�����p�{�HQ��#�p􃱟0oCqGs�zߒ�A���L�aq�f�f�>�f�F�94��Һ��	��<PΈ"M���Yҳi��hF��2m& qA�B�tה�y�]�؎�{�_��]vk���᫨��X���'��C�Y���}��З�1LJ� 
/;pB'��le-Ыf;b��v�$Ŋq�?Iq�AҜ�Dk�8�n2Ŵ/_|�5*C׌��+�A�G�e�t��t�,�z K�[gO���ҕ�8<�Y�w��m�{@�Z�m���+ߡa�g����N+aV^������"/���]���/ȴ��>��=�S�hԴņV���{J�O�����$C��1Q�?�cg���zC}�����lb�nK]���5q�&��#�=d�&�A���C�78W�cp���@�{���L`ЉR2�W@d�y�l�T���i��Hǃ��/��!�Y���}��U�p��T�Nr#��.�w�E�i!�d�
c�wVb4UC�+k�dج(m�?��#�(��1��,��DX����T[������w�M�*�]�"�x���$��6i��`�'�P�)L�A��=a U�l���K^"GeW��ɏTie��+K��N�0|�c��l���fu�����1��g�v�a��?��OQ|CU�@��� C��ϛ��d���/��<6F�^£Z��Gh��/<��z������c��y�x��b�Ƣ�p�a\��U�w"�E�;X��T_0�Q���̦�G��Mp/��.dG�5j�;{aTsT�Y�0�d��q&�W$�58�Y����u�,TQ�K��9�b'�S�w|x�I�����_��0�\F?�
���E��MQ��ۑ"�aEee�w5V������<�>Ԃrjv_��f;�;=����C&0�=\1�Շ�v+�����?�$bh)&�O5�޹�fL<R:����G0��6ȳ�C~�Q� "�@��t�}!�<^��2����
�ׇG&��x|O�G��7����vٝ-80�z�P7���T��Ϡ�ج5,l�v���.쨣Bj�oRJ� �����YV�q��7��
��T�i+�2=�pz �2����Oǿ��N������'%s���>�d�ܒ�0�<_3��N>�;H� 7MB�Y9����v��{py�B�C�0�s�ǬP���T)u�glV}�=0�'�?AKZ��EF���-gU+��O�B�H/�j�ĳb��0L"͸�	��Y�#j�>�n0���/�̋~gUEl��<=�>f�'�/#&��w�P�T����X�ɇj�NRI��-&�t��S���|�d5z����w�v8Q��vo�����ߕ��W/ɖ Q��b��!6tN�d��-�S����b�(_ Dy�*xÌx!�a=5#�2:������}���A*pe)>J7T�]Fg�H�.��z�fS|}^�:�q�x�bDN0��\��d�?��z�m�� �ӻ�y��x]�O��l:]Ԋ�Kr����g��e����T����8��RlE�J��A:9�[��x&�q�QY%WP�"����P�&r��m$�A�lm~`Z&n=\fw.M���]�D���g:��4��&>U�-���fY>+᜖M/�g�Q�I��1N� ��u�^%q��!y!y&�׮�<�A{�����ǭ��!��-�-�ڮ�����[e������k����m��	a�f4�܄4��N�C̙G�m#8&b����h��ˋ_H&���,�O]e�)*;�,����:��אQ�Z ���JV�z28%_r׫[Ʈ5u����%�X��̈�	F����Fy�@@��+K5��%r	ӄ���[�~Ż�W���Mx������u�Ȟ���|%�g����1&���:�O_����N Ine�� M��@Hh.[��Q,ߡ˼�!�)�!��3�Ҍ�TB�=T�c
j�C�3 y��'lYQ������*�'/>)A�6� @�th��V���c�Ф��S
��e�ۈGnG��<a�7�;�c_H�)B{}���k:�dPh�g��V��L���h���6T!m]�O;���S��ۈ�BR��y�6��;���C�`/ڂ'~֪ �!Ț&1�|u@}=��M5�fȆN��KЄ���F���J	�+n� ��7�ͧAn���(�?�x;P�fj��*���^|2C����	
�,���_���?-����w����=��������C�K���-���l� z!+zY���C�@��(J�sHb�|4/`�f*�82뇺�b?�-�Սn�a?P�lH�ނ����Uӎ6�_d9�1��!<�nӌ��E�:���]�՘k��+��.�"��¬҂�"�y�mԟw�!@�%˟�#�c����o<�
@5�1���{�Ld�)���M�O�E���	�Zzb�C��$�F���5<*Ŧ�d��;���DW��sM)�3v�KX����AՓ����ٌnܓ�8������ڋr� d��,�-���
t9 ;~O���*��	k�4�F���Ą������|��>A�1auE�v���[���N�:��!YaND&��?�h�]~�:<}jE�9R�u����wjD��B2>�B���Ð#�U{�]	!�%z�i1����1�������L �Ο	(��i�'�)�`X���fDT�4�ޑ�x\��M��U�� ��C��MiM���X��������L��cGm]4�u�6v��}��!Y�G|'P�����'�L��#ha����$�38��C���VQ�<ǅ�gV�f�"�z���݊����Ր�	��o\&#
DF��k9n>�kp{^�V��0�",���s��{Q3X0rMgR��hF�6�i�&@�x�󚎦3���82���s���T.}����"@��ĮZ4UlUuy��{�Fõ}�|�-$�}S{�8y&�(��?`m�H�y.��B�%ѿ�ڭ%�$��S�>QDD��Pαa�a}?��.�CMb���'? r�y�	pش"�U]��9��^�!�P�~i�S���N�ʼ�o>�~I:�X{͐T�N��j@(M٩ސ_�'%sGjY� C��F�(�u�|a������7�h7�Z^#QŽM4�M8R�YS�	��hb��=��w��;��R˙�WÌ-�DԊK���s_Up5���M��mClm{�vY\�^�B�͡<P�_v1I����5(�^\���i��K���m���Y�e��w�#ߛ�wF��G1QoX<o�s�y�yڳ�y��w�x��,2!�Փ��7��6֙��Z�-�%�d#�QN��0��H+r%�d�ju����*a���;qD�C�d6\ׁ�:�����N��6r����<�5��5&��JS~VM�J%e��{m�K:\7��s���W����gF�T�1������x�ֹ8ݱs�����Q^���m�YN-=�xZ�X5k�����l��ā���@ڰ�v���[�����*G8|�D�߽�����d0�dyP0�n��Wu���A�Bu=�����.��'Z�g�۾~���|�փy�
o����ϧ�!1��%5 ����WJB�m�(�=,3׿A�J��8���1�,BTx�<�^�CL��BqZ�2zђz���=���&�Mo�~yDf��v�*��E�wQ�C�&c<1*�jRN,��V��C�����h!%PP��>��m�7����RO"'��;�?�ox[B�\���J�y��'A/4�r�������z���K�H�e�3Uv�@��O�~ee��_���h8Ԣ�נ�M\��EU�l1ݱ���\}P�o5�cG�$M�[LV=�D�x�FH�U��z�����(��x���C�[��I�ڣ���g4L������v�5&����irF���>
*�rZ�m�h{�z/�#�0d))l�x����8�UJcJ�O��_�F�;',d�D
���z]�1+�]��6�$E�� ���-B�&c���������d^�=�-m�<F�dK���.�\�}���>�C�i��Kt�$�ȑ����x�4��<���!]R�!�—�N>ʃ��%����X�H_h)�h�2���"�d1�[��G�vQ�V^OHP/����2�A*���h�Iu���"�F����;y�Kz����V �Λ�������{����&u��{PMQM�	���\p�o���� w���m��0i-⣤B��K�F�(���q����ɹi���w{;�,� :7ŊdaMyAĵ4h�Ə�nۃ�y8�+X]��c(�m���Q�4D�	݁G��Ҋ�#�i��Z��V+s��(�EC��M"�����U?=�u祄��XY[��&�i�3(�%6�@$��������_�7/C�K}'���aķY@<E-b񸱗v$鴸B	e�M]��-�q�]���H[]�
�^L/'s#j;Ɵ]gD���VN���?i�d�]=�)L�O�}�#�?*'Y~'�1���#3���1Z �dn�M^Uֵ��ږ2�i���Ŏv�ӈ�U�_[��G@�Q��_k7��7#�na�׍���.�_E)t�dWRCa�<8D��ިgQ��;�iwR����)�%���<����|^vb H�V�.+���oc}>�&�4eJ:��\66:�C�x����X��Sl6`�դ�U���jЧhc��o��X'J�}�,�0Q��J�}Z���_$��Α����3�L ��P,�]
$�W��|��Fٿ�Y�A=5渨@�&:���ث�
��������/M?�/5<��B,vVUy#d)~wC�N}���<�S��[�l(y�J�*a�(�#�U�ځ��
�%Wޞ|�	�t-�C����9����/C_@��[�A\G�}@��L�+1��x삤E�j:e?!]u.�Uך1� *̖�]���d��{"����j�V��qnG�Cνf��\w�ж���$݅���.���t�H[F�N��pQE�nv�^]�x�Άw`�*>���n���E����^�����@�G�:MT�婢��ּ�����
J�T��P�5��A9��>�w�"��CIoQh鮽L�P8�3�6ZG>��n����GJӟ����H�<����[�+i�W��#��Y��A���u�Г#��D��xk��ML((L�ڄ��/��\���Mud�Շ@b1�P��>p.F��Ql�ح��u�\�@��u)��)���l4��q�_��o<{��"?ȃ��\����Y�,�6[��:u�\���=w8 3�D����1�EF�#�S",	M���3O��|��+ !��{Z�\$(�g�FGG(����ho��\)�G/�&��ms�����
�l/ͫǞ��|a��)4w��Ïٙ�YL��x��*o�}X/�^'u��Bu�ZȎ�~b��������y	����hϞל���YD�R�	�ma�ƃ�g&;� o�S���X�qͨǨ�t����x���޷�5�����E *�h���\lZi���QQ�$BH��U!*�(�E�ELqG�V�D�В���T���$�S��=���gf�����aR��U���}��~�J�/�����~.@4�"D��: �Eg����ams{9,Q��%A3�L�[�<x2I�X爳Kd��[��B*>��{s�9�2|oزph�R^��`�	���2�B��o��T���-V�qҒ+[̗���f�ٟ�w-�mﺘ�B;�"���L��:�4Ce{d�����Nv6kR7��z�g� 
���� l(F��F��cr�������YC��ǯP�Ӡ��D���*3�@$\����Ӳ�'v�ޯ��ߚ�B0�m�PFJ/�*$O^�5$��hҿ�A�0ʹ2f7�.������c=f�;�������3��mq�y;����5@*}V��>��M�jK<���}b���Hm�wҁ���U����&T�+v�?�CmCU�T6�L�TR1
3��be;���F[D��wK#��1a(���v�FZ�nM�x�=���!/�kvm�^z?c����E���Az2�@��2��G��mH��7�\��5	)�>1hL�f_Cn�j"T�����o�u�Y���b�X�+'�L�#��0����#�Y$�z)�5�Q>��"0E[��D��N+I���6l�_���Z	��47,��rTYU#�0M5�=��X��P�����y����w���W�����y�Ozߍ|C��N��E$M&G���:E��`m�c�[80��BK�>��*�?y�n���*�������Mv	(ڰR�_j���<�����(�[�_N����O��J1��݊�H2�p?�K�F�[/*�x�0�t����}�'�F4��N��$M̼{��^�X��ø���7�0A-3�0�{�M��V �y+��?|�n�����FZ�c�Gp
6�5S#�!uG7.��%�zs�yPUT�uSN�5;�����+�?C��.��ZNj[���'�!!#��$fPI|-z�>�|��;���MU�us�WnY����$���U���&�*�+L�W��\��e��"�ot>t�p-�f�a�v-Ix40f��.D �7���BU�*�ͅ�E��3��K[�Y�V�T���u�5J�"��$:#V��J ���tǀ�.u%>g!U���"��V��	CÕ<^��buz��LG����1�w�,!����+���$��:��Xz�<�Uq����\>����ױ7���sI8�'d�a�֢���?m/���[�S���S����R�%��n��O�1�9r+J��Bp�n��*�{3Sr(-����0F�;�_�0����m�Y�ƛ�&OֳYQ;T?#�Ү�)�Z����G�1���5����& n�E��K��J�>X���?��Goth���v�j]���N�"����l�]�e�m[@]��S"X��*� v|�"�p�:���-=�у��olF�f����g���a�����`J3>!�V�B��ܸ]��]�_t�ɾ�/H!�J�7岧-A�JD�=�~I�g�Ȭ
�pWO�����rJA��K�u%_�C<��wج����:P���^{�^Y�O��������a>d43h�a_��&s=����}���.\���<����R�'?�Z�� �(�"�b=G�U�C��#�l��Y�F�hD��D�ho��>x���O�p�H�̩"r�6H��7��~�v�j>LA��z����FV�D�x%�����s��0`v>���HV�p�U�OO��]Wb�F���͒.�Q���

"$=@_qV�����5�_'���KC�.kܴ�˦(a�� �*��F	��4t���l��L�C����w0:���
cv�[����~�������"B����`Yx����^�K�vO7��[�V���f�WNo,�o��s����~?�����-�J
���^ҵzn�~^_W��`�@s���Ɉ4'+zMvʘ��/�T_bR��PZ(=�"�A5�&�|�W�M3��[�xO����qK�[(��ާ���N��{�A[=[�C��'������16�h����:$��9��2����k�8�n#U���'����z��`[��J4R���om�tB�5�s<��$�Ҷ݃n�<��WNZ0N��ȜJ\
g'�Bs��o�I��d敁:���4�ۂi��cٷp���LB�QyK���¾&1�͖�����3�C�8Q�y�ʗrm
��_!�}����_�߰>�k�8�̆�:~�֮�e��a�߲�j�+��#�5�E9c;�.��
X�����V�H����I��{��b���+ʑb�zJ<}���HX��w��~�	fǳ�Z�$��C��q��ъ��=c���m��f�l*��$�h��U�xnI�iP��h ���Ui������pN~U;X�RE��G$�MmI���*eۓjc�1O{,໐�">fs۴k/$VxǢ1�}VI�#Vwp�.�e�/l\�r梎�-�=̾"��[�V$���.�4s����,����=>��Fs���X{��-/�y3S��{� x'��(e��Dҏ�yN/Ū�uum�ں��ı��jE�a���$�j]�?�S�;1i�������Ͷ@��O�jy���~@�Ť��w�����Ձ�'�]5-R�CI���Er���1�e�>q��
��7����Ԛ8��N��@�rQv
��*���)�Sت=�d�>i;���w����T��0�4@rM��1��Hs�9���O5S.��������+�����Eo1_)'�T
ddOޘ��g�2t�p��X�g*;/Ԛ��x��l����[̯�͏����Sf�v��4�T^�rg�]�m`P��0��D[9�<�P@�	+��Y��������>�Li�9#fA�l������P"]�����L�ݶ�����ʼ2v'Dݥ5B4Vn7l��ڕ����c��A���	�����)��� ,U�DK�k�\�w!l}��Hkb�2�;f�iK�_���9��f��ūlF]��S���IUn�y��yK�-��*'��z�+_��Û+
�iovK^}*8��]��@���2��
��+%e!��U{�G�p�`7ռ6!%��k~G#��o<�^�L�������0�A�.��/��5��q��lK���]�������sF=B��+1��Y*v���mr��{��`�tͥ+gw9��l�uv3͡`�Lzq&�1m%�pP���+���{C��V��dy[]����ÝcFڤnY��\����b6n@��Z�<ڳhp����z��?��� �+���H���|�h����[^�q�};s�����sE��a�~��P���p����'��������*!d
�1�N߄�D̕^5�9ѣR��<Q�ǋ��݊���dtղ��!B�s�Znh�կ"­<�}�	�
dj+��}p$��j�M�XA�;�I�.F?��@���:�Gv*���V=d/?u��+�Z�l:�[Į��ؖ�d0����p���� *Σ��a�u_b-��C]}��4�H�(�h	!^�)����kzso���ek�x	��1yK.����E�07��f�	��2�
�G��lg�������C�2���7�R��>+�sf]g!�����j�����"y�O��FL5�B"wU �p^b��_�w��7��S�3��oo�p:E^�A-����H�Vk���{���ȃ<�`	�Z������͓��2}��:T50%�k�ԉa
�Ә�����^��^m䒘٭�`�l>#���l�P�8m��6p��-j�޿k�_&/�I"U��E:�
���8���k��U`��f<�;�d-�F��1P��J�(U��{YAeH*R��WeX*5)
���������a��U����0���)3[z-�k�����V�+_��ZI;��t��q�{����B0�����_٪r_>��"�{4@���_1��������M��3O0�#C��F7Pm�/��	oܝ�9�V���L�h"�ϣ��v��<����:��:��؅[;0�w1��{����1��}g�Я&���S;����*���-�'/����Ѯ�Ո٣���< ,�^�Ù�B)���NQn�����ǣk�E2�o�E��K��r��dS�B��c���~����!85�åD���&G�ľ;I��o��|�neN�9c�֭>�ER��*W���/�1�=D�ܼ��0�x���B#:����~���o%kH�E�ڭ`�u�^���{�5 �p�OPeܐGj�^D����Xy+����A�����6J[�}x������_���*r���ؒ��I��#�C\�O�T�H����Rm�
�n�0ts7G�,;0���u���(=���'}�qqu2�:��z)i��~rN7?�j�WR���>�[�}���B�����ӷ^��=�[H7�#4V��\��Y,:�{��Š��Mn�'}��ac5��S~��?%�u��˧�%�?�?m�ݥH�T��f�rA�0�jʠD�.`i��?*@m*&�4�|�E,jkC���^���p��:�Y�+��Z�us�Hs"e�b�������&����O����b�����	_��8�qB�{���w�s���t8�h@���"0Wi�xN%��	��~,�%8|����{@Se䊺1�0���£W˦�L����k�C��>c�`�}�~���zk��ҝ��ԦQin,�U���`|x��.�)��&���[�m������V����pK�ه�w!S�%A�Ս��i�`)��j^ڍ�e�^���Q�.�o"P/��G�.V}��,� T=ʃmZ�p����<��!�{[������t{�vʢ<�Z��R�SQ�OO���{ �H���/�=�y��k���b�jQ?��zE��W��]����!��-;�NL�8!��n�WL~��8�f`��r0���Vj7`���:K��m�wr�������r�_�~����3�B� �O� T[a��!4�bg����S��d�홄��MtC����5�G�����b&;�"th:SJ� ��[:�E]QZF�gg����.�]#vv���޸^B%^f�B��z�8�l_���2�&�n���x���>�����tT�"����u<*���}`K��kԍ	�P�kס�P��01E�搝�U�:���&7Ȣ�s��2��Ӝ�K��Crv�eh}0�U��SZ�ǭM������O�R�|x�-9����o.��αG�@ݠ�<9�X�S�/�	�	������-�t���i�(�-�,�^����#t��Q��G�:'/Y�_,��6�gH�ã������D �(�*�;6O&��K
�7fߺ ��ç�ƨs��l�_��^�n��D��-���Sک<���2ah�g�(z]n���~#S��n���~R|�,��pg�*d��b)En�M(�?������A������*��^�4��d���\���n����f�)q#�Y�A���u����}dV���B6�@d��-o�Q�(�"L愚*$|h=��H�~",~j��`"�>
l�z_��)�1V�����OvT[��,aw�dV��⻲��)vf֍8+���r�E�|UVo�C|'N��N��p��^�� g�re�@w�ѬRj�.�'Ύ�Zc�Z��[i���]�*r����(��������j��~�#��5����n��U��{�����%z��pO�n� �U79����R�E",SoG*�v���ͥ��tu=o}d����­��>9v�9� ��X�}����/��X�$�L�na��c�@ (N�O��K8Ap������C�i)�6�������w�b(R���`�5U��}��$�i�r\|e��Ri�������$ފ��!�ʘ�k��8����V��
I�Sr�=Q���<�g	�5�R��ߊ^�ŷT�@�n����c�����JBB��o�ԭboI�P�Qm+[Y��x��+#,���{��ꮬP� .ٚ�<���S��	W :�[�"����V�t@�~fw3$Z�\�3�-���lu +� 	�)X���[i���-	���2v	ɖ�b���6����� �O�R�y�h��Ub������e�1�`��A�hfVF�3��=��t�б{��*��ӊ�{G^;���U�"ĸ&�����$<�"P@��ˌTj�����y����Y>~vT�Β'�1~����Q��9�b��cm�"\}�i�r��V$�
BkN��!�ec�83�$ �ٙ��u!�/rU.��I��o�him�Xf/$W��tE�1����OMy�,<ߎ���X�@n�ɜ�W����^CU�2?��і�m�P�f������o:F[
G���p�`��Z-1@_�VUuq,x�;���I�J��*/�$�)�S��sc+x���U���ő�����&&b���K��r&�c�� R�`�P�\)�v*7I��E薃��C����5���U�~E�)�@a���Ai����Ҫ�2;稦��"	q'=� �>u�����@V��_�2�k�/t�=�)����;AXD\�i�_����h[��Qm��L�q[&��l��dX^����Y�����2���
�O����#v�ݽ���0���_�h�C��VZ+�|�0�uj�7�}SN�&J7��V5������Ƭ������E�Պ��;v�5�#�S���[7���%Y��_W9[���9�,v����E�����o#�J����x@?�r�/%O$�SF�ع'�	lF��-�˙��f�~�`�f˟;9`c���$�;�)�,��Br���eQ-[r���d�|Gm��ѥ2���� Wlf��E�YO����ï<�4�U��D���� �w��F$4x�1�HzT�=&?��}4[��ηx�7j�śLA&;�tP$p��o�槳�!�#�g��b�
�_̓>�b*e�c<��3ŀ����eFj��HC�>�2t@�`�?�il�y�U�ܪ�����sE��y(�iO3��8030|*V_/A;
J`�R�n�-R�:J�ev0$�N�|�0u��O^{g�ܡ�)vؾ�(��Wx�y^������gwx�sT�!�R��}#�� �`O~�j�f����`��s�>i6��)"�8W=�u�g�j~�#�~�m���.�?#�?ڷ�aw<��΍dL�BjNgaa��s�7*>����M�)h20}��6���*�B���AM�Gr���Z*7}��Y��Q\�/H��F)��bd�p�$5� ��֖�����a��Q�p':+{���)8�!lP�Ä�4���~
�N���䑖ܽ�}���,~]�J���T�[z�y�cx}��4�L�!P����`���V�)3�j���r�@� [�v��Gb@ռ��`u>A�?�Z����t���5"�#�9�_��)�5��G���W���m���SR����&u�x���������c,Z�o���$�Iw ����#�D�I6���5X�������������R�wЍ������VW�r3����z)�jЦW,��m�艾n���d���l�:��[�Zwǒ%f�IN�J)�YeԐ���M�M�[ȝ�@?$�4hGH����>Z�C��÷0M�N����P_��{�a���p��-RY�F��.�h���_
��gO5	`�;��/�ܥj����֋���=u�nL[8�&�S��&�);,����*+=�P�0;t��1���l&$ES�o)�ga����l���=U�i���l�D��n�&<3��;'#s�Յ��c��cC��XX�=(�ȸ��;%�YJ��i��fֵy�+�g���˺�k��˞��#[�&��Hl�xǐ�\-��Pԃ�Fr3�w��ry��7�pDsx�$"><LZF�SB�V"Vͨ#.I��g���G?R�r��s�7�eJ9{���P�� �Bza��O��v`{l=�h��ٯ�o�+�7�btl�@���.� ��@�;n�V�v^nSO1�� ����`*�$��nޮ�������s��{E�1�����ú��7pص!�!�w(�!>T����	;�y�pt��T�ﶋ�l�f]֋��_H���%FE�i�'Y@�W� lt>��S�5 �)&��$ڧ
���x"O�  �]��W��S�[@�-aͯ��U�B�Ąs�o#s�M�Y��j~�l�l��x�|��N�����g[���Ӷ јnH���T��93x�f�;ݠE�9O������q6_���1�j���oW��w'V��q1
�C;#-lU���3C��@�(6G/Vȫ��v$��0ybi�b*�����P�79�yl�e�?�k����%�g��1#��: �:���:���xĻ��!�R펕쫕�4�yU��;O'����}��M��y/�"�� M���.��؆&d�λh�pbg���UL�T���+@������3b���H2�s�B��?��5����:�ww/�N%h{�<�9����#�t��R|V/vH�����1�� W�&O�O�����D��I"��T��o����%TF����t�+�1�4d@�	�~h>r@�z��
��޸�0oKd�<�b��[퇥���O������T��xb8�<U��ø���Z��һwT���N73�$�-$��*9�t�����.u�����+�n�Fu	��}-3�;�\\r��-?7���'���31(�L_f�D���_�����C����2'�k�.�\I�*�L1_��i��ށ����>/y����Y�X|`�Ձ=��6�z�ڭ��[��/<�ߺMq5?h�s���!���%���VPZ��4�~��ʹ�du���#'pA�����0x%N�7W���܄��r,_v�t�^j���-�+\$�����b�r5�Ѕn �
+~E5n�O�oj�G�^��SVf�Go��Y����UȨ�&��5�iN�� ��r��5�;�$ 9��3����pf�:WL�G���$�*��C[
W+�������J1�D�m;o�ɹ�bR�ɾ�q'3Yv��/ݼ{�����C�S_g���R��2S����b1}�	�͒7��?��y�Tʰ[�?�Q�ƩR9�V���GTRP���!�=�~
�R�*O�"g$R����q��G\{����$�>xp���jz
VV�!{�o��H���z��NG�h(?��S��"�n�m���ϻ�B(5�:'�!YMn芘ӹjVY���(�g�+��G�� {r�:���i�﹤fc3�� U�d����d�-�u�v,��]���r��A&.POl�	�S��{�
�8_�u�IV�u[F���2����TV��.$Zƭݭ.�nz(�T᳐{JMU��'b#r$�״F�� ����Q�OPZ��|@�`���Û�g�nu�퍱�|֥��6D���p>��"9^��o�q���*=�7�I����Y\L;N:�F���JV~�k�th�-UF��MYd�؄�u��i���V�M��>���j�9��T��c���ٝvJ��Q���]R��m��n\���c�l�s�f���D�ή�,�s�3}�\wa��<#�������"��*#+�O�Y����e�=�)*�Ij�S扶�G��a���iư_�{K2�U�,��sF{L~���l�(��n�M�d��"*\���_��6հ������(<r-t=�#X6Pm�x����*�^�@��sҖX�i ��� 7r7-'����L����Q�7RM�`�x_��#1�ĕ�m$}���b'��BNyqUa�g	��߻LO��Ӷ�b�ɫ��9%�2	C'W�=�����&�;�Ⰳ[&$,�]�I\���\aT��j[����g	��nǴ���r��F�w�2��G�y��3�h�|#j�����R6�>���SNN�IBb-)Ht����V����)�-?��\L�Tr�j>�ӄ���P���_uH.�u#JYק���N�0y�I4G�v�v����%�s�e��ٙ���/h�0F�@HN"��ى�=z6އ�m)cI<{b1י<�a8*����}�X�U�p��p~*������A��9��E��N^��wG���rfS�,�mp���<�G�Tj1��������C)�s��
��.zE��-qșpT�Rߩ5Vn��@���Y%�j�������u��b�k�ا8����w�Ou�.�	|��L�R��ٕx��`��x�����,��2u��vY�h7�g�k��ɨ�b��Q� e�vrc	B�c����%�>�����pB=j�f���'We,��x�+��c�N��]�҉��c(I���v�&�s�&gtV���!�؇s�m�W�U_�f6pj՗!I�8b�;'z��X��#�e7����=OL������~�����a��(R��R��7���Ň�~^1��X�9o��$���NN�yޥZ�lǆES�N�]b�y�B���\9ߜlD�#Z��PO�[rKV�H/���`�Jx�n�� �<���Ì�;;���\^���ȕ�'KS����f�}~<�3C6^﷛!<�8&���SP����{C�B�G�]އ���Y�%V}���D�&��W]�څ� ��į�NV�.����5??U�x�'�G=]%�uA�������F\�u3g_�d��(����Gh:�3�/���HĽ�g��Շ�[r�U�3��?�
�z��S�Cbr��"���yL�&�oBD�ӽ�$��0��|��!�%��ߟ����I��e\������B�Nv)�Ю����į�|(lۉхs��>�H���:��:~A�[��0�4��z�Z냾17㡿���f�U�azgY?�]п��&�Y��Eۚ"1��:*���r�Z���W��"���|5��T-�Fe����g�D���#h� ������+�?Y#[�D��)�EH��������Vle5-�kμ�"HM�U:F�HD|_��?�a�ۭ2�t��{W��!=��d��=�_�|3���cttZ����Vw�<bWG�-ts*Mϭ�i[-�~J\�qn'�E� _t�}��}�	��P���ֶ�g��#񪕝���S�_��-wg7g���3�`�3E<����b"�:ہL*�5s������j����~7~}��v���I�z�=$���C���1%e	��b;3��|�>k$�iL�������0硸Om�{�gc�LnL�����IK��h�&E�Z�)��is%���h��������:�"���)�Tn�P����e���=�L�T-�/(+���<�K�@2��.������� D�\��򆶕��B״�bj�����H���6g� h�-$կ�ol���z������L�}馻,�`pD�Ĩ�A�� �$����@����^^7UU1�}���>Q*�U��͠�0
T/���tR�\�_u�O�j"�(�=NV���������;��<�buEI��$Q?{��ꦊ����]��`3��ū2	5�Ns�]59R���f~�Tg1=����A�������*�{�~�L����A�5y�"̊��,_�����d��[避��Crl�d�h�'پ��$�\������$���+����++�,�-�5C�I3*Wu*�C�cF����UƔy�o�x���^a7�o��c#�/�-��R�B���eR����L交z�X���I�A��WxscL�8�$2��Ԓ���E֗{�����U
Rs������C|�������a>̮c��ꓝ���H��
s"�f��e����2Ő��ߟ�[џX�
�?}�XJ�{Y�\}	�`&w��z� �\�}���x9������#{�A��ڄ�c������CbZ�����>��Ɔf#A�s5�E`��P��}�g���|_o�L�^���:-T�F��U_!9�eMy���Í
��b	�k�'�)�.������e��~����Vn�d��H�k��e���x1�`���0�$�!.��C�#IBzM�}�-/�,���6�<�0���Zm�5yޯB�GV0[�h~��8�0?����i��s��p���]z��3�y��e��t���n�X��z��w�/��7�G7Yw��p�`�|;����^E�ryV /��%��hNrA�ኣ�+=M(�t:s��=#�
�A��8Ϣ̼S�O�rFfrV)ƿ������q|�ζ����	���Vqb�J��'�b����W�	��+��ͨ��^H
�2�P��~��<�����|t[6侩:+%Iyem�}ӣp9�Ā�O���R?�o�ϟ&ϥt�z�_,^})N������Rۜ�v��&��G�\��THl6�MGjO�z4g�����Ώ��Z�-nm ��|�>�3Rv�s�/�Z��ˬ+Z�G7-�p�J[i�:�.$e��|�!V?��������\|<]~ðm��c<=���_�����W�w,���T�������F�<��JOp���>�-���{<�ٳ4�|r 0Y'���:8�[�ê� �&�'�����MYH��4��J�j2+ʁu8�j$���Ťאq�����	Y����R�������Tq�r	���U.�/��T;T6,j�/�Ƈ�����lm�ւ��9�`E�$;Yek����}$����7G({��\�P��..�u��nHN���k�!��xҨ{���IY�3�љrRS�c���-e���}��(��r+b��D�-S9��4���1<�Xx���;�<���tsүN�bBJ�"����V2�`�i���J+��Tm���L� bR��d�~����m��{�uY����`4����G:�*W���&��l���ʌ�SO�~ɉ� 8��{�˽c2'�Ϫ&�qovM��S��P����8��1�"�|dWe��DU�2�E�-��ʳ�#��,�ޅ�6}ˏ8{���c����.����3�������	fD�������o��s�%�!/͛`ǘv?�AQ�x��\�$Lp����]6�c�,5�-+T�P�lT�6F�K;���N�Ȁ6����j�_c���w��	wDݭ{�8���(��{�t��5�`����c��az��.���sC�j�5�r�|�#=�镟��[�!t<��Q�~t�}��н�E��-d�	�7N�����P~���|��&t9���F&;��͏F|����'b�'��8a*�+���`�"r�bA*a&�Hm{��X��WF��l=[�LX�?AƋ�.(���$���E?<e��W,��,4����ֱo.�gi �|����%L��r(
�r��$�A&�EP���[���z�w�[��1�~}���m��hPqJ��I��Os"�^�#�S|���nbv����<�죅b��� 6�B��6c��0F��?�(?�{�r?MY�ozL]S���X��Ua�Wj�12�ѯG�Tk*�٪5b�,��L��C���C��yQ[��O�/�����dc:�t%vs��m��NCM?����������a�o��~��]��)i7�h!���p����`i��]�h��8}��]]H_Z��g,,�i�E��j 
r4"�0�5�Z��R /�����#�
9��7�y\�[�����Mkt�A1#'���p�ڨ?'�jļ�.�d�(P�d��ID����&6�)��Y�gs���]�8�B���t'9��%?r���m�5���]�����+�+�<%'�Pĭ)QV�]�хo#{܈�O�7X�Z��	NwnBV�q���Z��ʯ�E��ӷw���P��E�q�6r��7���*�̥-bǤR��<=#�V�[
�R=��^疭��Lh�w!���\�3���L���K/�̎�l.��3jc�r���mY��,�_�BlmޟO�,}����.Ǐ�#f��G�;��k�o7��Cn��7�Čw~S�ʎ)�GY��@�X�a��~�0dd�T<���حw���$tm3�$^�����ݼ�M\R�����鏪f��JA�@A�c��a���@�=n�o�B/�0\_�PJ&mBs�ɕ��w�U�#��ksO�yh3�l����˃w���XLv:g-ղ���8�D�ȍd��_�Z(|;j]�m]mM|0Q�E̬N�2#�t8]|�˼��|ħ3��|��K�k/�덧�x�p��xxs^�*I��@ݨ����'�\��5C3h���"h.���Q�S���]u]���ZgS?��Zֻ������ 뤪��[�#�n�$�a��xq�<�����-[��ܘ��3�N,h��UM��ߴ}ؗ�V������+�S�V��~�w�b�sSzӬaE��,�qc�\�o.U>U|S�Ȝ%T��8oF1��������8�h���۱z��UfE����'�\��~��ֲ��<��/y��"F�1;��G�`�@e�bBa�;�֬]�{��Ȝ!�iϹ��Ӳ~�"�Dp��Ý]�:nZ��d�П���cɸ�k"vrU�oI�����U�,z s��()�xg"�3p�<��<+`F���tS��p����Ɖ��:���\�y�nOm��U��v���6W>����q1��;�Sͳnt�/C���Tk_��`���nJ�퍳ꅂɈ%��C[�iS��86�&)���׽hkO4T���A�W��*-��[4[�+��E�ݙ|7�,�Aa|sR��08�F1M秳���N�����j�M5�B���������X�D\����y�[���׈�0Ic�dP�W�艄�T���Qa���6S?~�q��{��=n����m�����1���}.&��=���\�l ,,�JAq0�h��u�[���A첰T:�"�'%�I�/P��c')tSD$d"n���y�ZT���hd�?�#�T}5��C�B���LNFT��oW�9DJ��z��B�k7!i^�ɉ�1O7O������V2��r�؃��4�"P��7'�E+�[�f�P����ѿ�j����Y��NŚw�m3�1qY��,��.ͽ��c�:),"]��
S�-�'�\ߦ{���=v�\i�~}_�#}���p?�\� z�_��~��,x�@�~��%z�SR�@=[�R�z���oK/A~7��Li�"3�J��Emi$��Ee���B<����]��[���wLs��F���k�P�O4U�`�t'�Bjd?�Dn�:7���9���g1�2	]C�w*J�aeS�=<Ã`�������B�,:3���Yn���������O	ݖ�8ì�������_������n9�"�d$�6IX�Y��to�f4�߉?�y2���ޙC���5Y3�T���@��5�uŵ�p8��0M�XE��b\�'im�Z��Ν0!��o�|&�q���*�+�n�7`�ٛ��|b�w�&�l�]��U(� G?�UD����k�eTaI�a�'�S�W�*m(��{y�4��b}>\�J摪p�i�Y���H��G�	]/��ť���Zl'�wo���g9+U������GD[�QN³�ʃ���-C�����vB��i��h��(�1�@ޚ2:��v(ќw{��g�ҕ�gFZ�ǳ� u��<��5�Le`�'A:�0(4���O�nj����}3uBx�� �7�M��etl-�cZ��$�Z����"6\��a�����4�~BNI��z�_��޻���*;*.ݸ�\�O]4���?y@�D2�>݂�,m����i�����xY���@'V��T+�H�����ƘVW�f?Ʌ�^4�-�Tf*F��K�����5�P��6�[?�޸�(��7qbkբ~������	1fSs(�8'�2)g9�n7�'q��m3��NN�::m����W_Sǀ.�m�:ĭ�˒ܒ�G��}p���,n�H~�r�4�$W1�X�e)����"7��UL�~M��s*�;�{��k~��T�id����+���v�C��̲T��U!����Ԝ��rK�^md��o9;�4t��I�>ҿ����	Z4� h�'�:�w�|���Ҭ��{¾�	��&�v�o�B��C٬�G���A��_C�?z�i��.D`jk�c����%C���oq?�l󀘪z5�-����D7�����m2Җ{q[�B�(!��/)�	=�-d)��;�t���)�P����Ӌm̫)!��3���K�.��w�'<���<��C���R_*7�qiD�T~� %o&�����:�>A����U���Pp:���&�w��n�Wn>��>�Җdq-�&��4@��4�b',s��[��O��@���B���^��e�B�1�!�w�F4"�ֵ4�O����l�	"����b�_DI'��$cjD���TFe��\��M���te��-��V'L4���9b1�U��6�Q4��P@D<#�_���TRi�+���]H<t���~^*j��Q������
��}�����n����&�x^�6c�]�,���d�\{@[$��p��y�RbE;"�����6VY?��ݽ�̤�j ��]�BtfH��	�k�r�,$��:�bf��������־���\$M��ط�'ʥԧ�H�r��nǳ����:m.���/�D�\R%#���2,�5�@rN]��l�ɡZ��
�'/;x�>W+ꋧ|Gh��@&̬Ǧ-o8�Ks +J_X���@�1&_�H������*ںČ��2��W@��o	�U����jo}`�҄޾��%���y;��M���
]���u1�:D� h^�v�r:�����e}��[�LJg�>C�e;g� gF��`��Mul���όo��tW�R���H��S.h Qm3��2.��xA-t՚dl�P�ӻ������}�P������t�T=^�w���p��'�(b���a2h����p>o��k�c���m����q!�J�!u!��j�P�?��̭Z���
]�b�������Z����?���W{��ĕ�GS�����N}AW�Hu�1"HJ���j�F��b\�-TB��V-P�#���	����+�r 
a!��_C2�@&�xzvk�{v������33g���|�~���~��E�cp}�`� ��]�����ڞ`����o���� ��Q��j�V0�>����i�z��uܹ�,<��0# ӎ�<��>W(hlƄ���(�T���X�Ӿ�kM��~rSh0m��QZ�;H�=���+K�wNx���\xϐ(���-�m��`+�g���>Ҙ>�P֢IT�m�a�{{oኡ������$@g����`1�q�'�v���W��z>"6b�S+�-N�.�6�:ٜ������:�	��π�Z�����<����BN��*�.R�Tr�ݽ�<��D��ӟ����q��A��k��b�@�c# ��O�<l]��$|=ZUu�|�Y�A��Hu#GT/�PYs����QF�0�6��S��`܈t�rg������{������t;I�v�2���8���?6 ���)�ǒ���E�B21��8e�w���&ʕq%�]e�c�	��?ހ��5U��]�VD�u���R������H��aP��;�
��	ƜB≷kB`���i��!�헔#0�Q�5-�]�d���\�e��O�G��w.jR�_T��h�*|�dh�J#���`���WQ������B��T��muf��?��X��JM�FB�y�3�����/�XpT$�:�k�x�B�o���o8~$���l��M�D��F%o/1qs��LH({^�f(͘�Tt�1w�Cέ=�ó�\p� _��9�����+����&a��]�zJX�'}>!�6a)N��m�,�j���&uL�
Z�
#p�����^��S�l#p����j�Rr�nh�ё�l����:�/�P���x"��i�5��6k�����>�eG\��֤�}^f���#Vx�.��D��B]�m���HZ��:u8(�.Q�Fu����ib�s�wj��jXm��C�䓇�C�d�)���p����;�~ީ>��d�W�IkdUVT}���~�Č��<+��K},π��d��~S�;����aҩ�1��V��%�Z$l��cZ��+?�0����?��U'���Aw��C-���p|�X����w�k��N��9�A��-�Ŵ1fj���7�1�,n�>X�G�V��A�F �r�\����HL��-o�M%��qm�����K�!ZlfVzc�����%9���v?U�_F�
�[�
/���J�b!�-&vT�����v�d�"n�/����{z�^,�<F(����~�	�W3�M�F�f��`��Q��?��?�S)^�S�&���UZ\���ǭ,��JO��״����_P��:
wZ��FC߀;Hc���Hq+�X�2�2�8��8�P8�Wx-e��@���#�X�����"�R8S�;kߟOO��,X�]MF�k�o>��$a���%'B�~m,ٵ��>��f�*?g��k��t�����!���Frv:nN�}i>Y��o-���sS�_��`��$e�0�Cd���߄�=����'v� !&)bǏ�h����"���ߪ2ط�.����j�k����0uQ뙫n�k��%����&9��K��R�����/w��k�{,[^T��Y�z�_x1#���+8{g?Bz�����Ж�ԉmKʛ!�>��3��{��5�C�&�(��d`d�1_�y�.r���ȟ]+�#j�%�o��`�zH��Lb5�z�/m���Յ�~ܵȽux��P�I|���^�k���|��[��͞��Y�*���.�����
���_�ֿJ;�C*�>z���>��[����tx�/&i?u�o��5���@�Q�wPK   -�eT�k�X!  �     jsons/user_defined.json��ێ�0�_e�k@>b�����^���[�RU��k(���(�^;i��`	���|��̿ݮ�`�V6�
����/ٴ�2� F0B�N�g.�����Ň���{DxmC�۪�������x� ��9!0��0#H��fy
C%�PT)���场�^�}�Z�y���$�E�G���G?�ͫ��7��=0��Z�u���V�}=�xDq"�{9{���FM(�'ĩ��?{+����F�����Z픾ץ�b�E�� 1%	a��}c��Uc�ϯZ��t	������W�*-�9p<�}�d.|�t��ЗΦ���/:�Oѩ/�Oѹoe�=�'C:_�F�/X4Ҭ|����>�援����h�k�r3��-_n�������b4Ҹ���7�e�xZ�Ϻ�k�`o5U-�NW���yenܣN��V�r��e��1�xQda*)'q����+EDy�f^`>��5/�aD=v���"PHc�^ �$�T0`�������^ �*���Ŕ�
[L�p���t�	^L����}�(�݆���7PK
   -�eTv��#  h�                   cirkitFile.jsonPK
   �beT��/J|�  v�  /             P  images/265b7ddb-a887-4736-b161-f7ff4501cdab.pngPK
   ǕeT&č  ��  /             �  images/dc330bba-b31f-438e-bca0-f858f4ffe113.jpgPK
   -�eT�k�X!  �               *A jsons/user_defined.jsonPK      <  �C   