PK   ��eT"�e�  ]�     cirkitFile.json�]�r�6~�)�r]�%H�6�{�C2SI*{�]*�Ǭ�%/E����ڗ�gZ��-�$Ė��j�͟F�����n4�/�J6�Y���쳩��j9��|:��U�������\����S��'�_�yT��h�l��Z�e=#����<byB"�$�tgQ�cV�(+��\��M_ݜ��C�M��(e���H3��r`�H�1��6츈	�Mu4'if;6$�\�h��,���Y:AH�<R�z��5�t�xz5&��*�Z""�3YJ�,#4Һ�q�d�e����0Pc� �o��#���)Fj6BjBFj���c���c��#u��Z!�����bԅ�:9��A�2n\�O�z��`V��t'0]�V8����vY���\E)Q4�Ĝe��y�S��)Pר����FJB"&e��I��IQ�x�v4C*ܷ`���)�g��<�D%4��hZ�Ώ���&�9E�-�3ݦHc�f4Jsn.�y���G&�k����>�k��y�������60�9�-��с�S\s�IA�k����7>�Q��A��*�W��}�	8�1å<]�`�.�����'b��5��@�!��'��#S���Ԅ=9b��ʒW{�}AЩ�t�{j�+���.�__���j���Y��w��Ac�q)
$��B	�=A%4�9��I3L��B�paA��ы�E�ᢂpI�pI��8�p|"���6Ȃ�6|�4\�_dF6 6�(��#���"�`R���p!�]�1lv��2T:nD��x�8�����u	b�2j�Q�q�@��O�p�4<;�]h�u����q� �������0*	�e/�e/���Ʉ���%�'��B��u�k�uʗfSWz�t��\X.|��)�s��)�s	����%�E�ᒆA] ��A/_�4�i�0��;�x.��;�x.ad0�)?�]�S��2��S��2��S��2��S��2��S��2��S��2��S�粯�/��u�'����m��SY���qag@>�N���M5��A��b|�)f�.��gpY����)Tϸ�5�gL�Q�z�Ԯ
TϘ-G�������ג{�3��\�|>=�3��AŔ5��7Lט��^�aj����R�U�j3T��S7��
��@��	b0�B�w�zî��Q���P�w��OzPI&�Eum���2��6��|(��B�]Pt�z�Ip���l@C��\"R���� �&� ��	/ 2����� c*� ���lv a�M h�uT���[x	�a�Q	.}�A�Q.���d������ ���o�����nI����0��F�p���El����P�2�#jS�*ߔ˗
���UQL^�7e�-�!�������;�gz�p/�e7�;��a�֝�N�e�e�²K²K�s^��ᇊ��ji�(�xfЁ��I�Ё��~������������.n���p��g��7b��Wp�#[�ZG�Ӂ�1���:�x�<�ֱ#�ǰ��a�W?��Z��i;�ZG v�E�v+�~��,z�2�;��!wl�܅#����#��}��9
μ:�5�L�,!��Ӊ���5rzs�νh��RGIi�A�&R���:���,��aױm ����1%�!�j�G  B����M����f�wH:��}-[�_�Q���x��׾�A<��8`���>拏ػ��0	TԂI-`���&C�I`bL�ߟվ�]�*��裾��,�{��Ob"�����+��ʳ���p&������˦�ܒڽ���s�h�Ԟ[2����ܤ���-ڿŶ�X�����[b{K�o��-ٿoo��[j{K�o%�[�s��b1�WF��\y^��-�u��gNHZ(ʣ�0v�ĊEs��$.�Zǚ)2����~�6vU�:TD"fJ]��?b�0E�x��}����Z�k_�K�գ��Ҹx�}a�.���H�v%]�Bn�9e�4�0��[�.�s��E��T�$�"�Ʃ��H�Y߂qB�ƅ��z��m@�t��J+�n�l�����>ˍՈ8Pɔ3r7���P{b{��϶C����;����Yֿԛ�\����6&�\q;ޣ���*���t+��J����)��:Lc�������C�2�&�#�D�[��Ԝwu�� :��U�4N���r��eb����1��d�X���6�Nz�[���?k9o����V��,�gr��=�k�q��t�Y�u]��OVwK�������^l���ٮͲ��nb�����˿Z���B/���\��r]���Ze��)+cG��S�B�A/7���Me�c�����K��jS���/�kc�/�!�#��9��"�np�+AOY;m�>�U>7l��;ѵ5q�RvJ��Jj��ʺ��	 ��B�9�6�k�7ŭ%S�x�4�?�'�*���v
gDELL[ƭI��yĩ��̩�⌫��y�ͳ�̋�i% 0`�з�=�*qB�<v�U�r@������	�s F�g�lWG,l@�?0l���&N�Xx�����4�Mn���	�p��6��I��j�l��}����Z���g��S�g��8��q�Z�-��#8�Ϥ��{�^���ͺl�oo8�����e8���0��w7���Og��tG�i_�?��'�7E����ij#(�IS�2�����d��WO˝T;��P�{��G��u��rŚK䊶��昹_�)�ޅ���������T�>�~��|}T�.힔B�0r��?D:��՞��2%����<"¨HJ-#Cya�,ɤ�B�oYg�z��[���ҥ;V�gU��O���N%��^���D,���͂�T���{�X\��7��{S~�w��%�v�-�߻-��g�6duvo�^�-+S��V���W4~��N�/��N�o���|;��Z����c�|�7�^���03��(+�f_ë�O������{@�W������ٗ��ۉKo}(>��4���]��q�R<3��3;��t�(�CD4U�S5�������z;�jw����!�CA���F����N�A����.��O�d�Q}[��?A�K��� Q	:Lձ=�a��k���<	<'�
<�k��d����P�*�aht�|3h�ᠡC#
ɠ��s �Acp�4d8hā�!�B# �@�H�C�/204DPh��0h �<�㥠��AC�
�́d���R������6��@#b�c$�!h���F���F�𖅀��AH�A�/0S$(4^����p��7�@2��� �w�$�q�ho����.S�	${ü�U�7��	��)4�ŗ/�IH�FuX��h�훀^p:�b�E����;u���i���[�j8WqX� ��� ���@�����	��q�t'�3L��K5��ځ��>F@` _/|+d�"�y��@��'�AǨ�-h�^L�"�|����Y�.���2N1/�e� �zݰH�ǂ�a ��� �+��L�	�[t^e[����@y�D�pO����!�3`v����:A�`���$mq�X�S���G�ѧ�F���C�!�q�~�	��ƫ6̚��Ayw�`8�Trp��k`T�=�\mb 4`_;�v�O�-4^����<��RŃ�����T��ʣ �SyjF��}�" �N��9A�` zU	O7BI�mK�J�F�j�M���PBBㄺ�d�W�u�O���Ry��PT�^�)�ŏ�6U��ɵ���9)�m��r�?����a�D��:��?PK   ѕeTד���l  V�  /   images/96360f2e-15f0-4a95-ae8d-a24fd3f977b3.jpg�X���6���
һ�"�נH�Mz�jPD�((�)Mz/RE6�I��KB�/��>��Sޯ���_������<��=e͚{M��3\�����@ �1�`����6 ��� �  �l�:6c�p�i�����
$�k�
�.��~-�n0`�+	6� �L��y!r!r!r!���������;������������� � ����� �������d)!!!)a)Q6A	)1)a  �~� ��@����~���1�~-s������:��  ���=��;�I���݀��q�H�;ӹ$��wL�B.�B.�B.��n�;��y��&!�2�`�@�T@��>�dz
@AA �+(�a9@ ����`# ��4@1��F��+�e38���
%������[3�-��W�w�� �	�	�`�K�D$T�$��$��Wȩ�XY����8��خ�bgb��qK@PDD��KRVBH�OXD�g%�K�.��Б��	]e�*��,���۲)\�U ��K´��V�~������O &�DD�-Py�c\\<\||<lgA��<
|ʫ��	�<4_s�z�A�~���� �C����%"Z:z��\�7n����KHJ)�UTRVQ���HGWO������������������"�e諰��7	�Io�%gfe�����TV^QYU]S[������������������Ʌť�+�k�����ãc����~a�&�w��������_ �(��
P�~6w�rM�!՝،�/�؅���n�D4"���]��g�s{��ճ?:��~M$�X%���  �qa��P��}��5D�{�F�8ui�f�dD��x�X��˹ky�_:�m3�����v3"����fڎ���,� �{�S<{Rl� ��bs.�x��@�%�c�yMbp��4�_�a<�����l�'�TD����蹘�?ؚ��1�E�_� ��0 ��8ʦ��܎F(_�V����y����,&�4���%��~+��/�mܝ$�э�C��i� v ��q��"���N�	�F�|�N��QΚ(��;e�İqs5Ԕ���K����[)-�c�]�E��+����NΑ�C~<~Dčsi��#���ؗk-��=��{×�&���z#� ڍ�@��tP�`�5�8�6��Ls���T~��j�rO�d����i�S�}R��X]d�ޒ��w�Kk��ɶj*7�]�����T���\#�}��sݫ"�58�5���(�6�t�u���s���ٯ�ߩW!��TaXw={���p]H�tXќ]/U$=���uW��I�l�|~���7�=��n�R4ۤ^2�i���%
������MH��?�Du���SF�����k���?(?I����a��u��$]�jj�4TY��	a�E*_�gF�{���?c��S�UY�t��l���ᢤ�<C�AǖU�K⧡��,{���Z�W���9)�y�+�r�5N_�<5uSR�'trㄿl��t������h8��}�'�d9��B"�?D������pd����S���P�2�
�
�=�'DI�^���O.���z�|���F��d����3�B^���wp~Q����\�#.�x4V��YSg6�h߀�*������t�;��C���r�j��ԝej�=��p��; �S?�=?D[d�M6�6n���y�Tܡ΂E�k��4SN���W�Vo��p1<d��	~7���d�L���r��HK �i���-}����Ѿ-���JnM�g#�g8��6rc�Ҽ,߄����Ӈ� �a�6g�r����'#�ܳ�܃�g ��G+�b�M�<���2���G�rc�GZ��Ʃ�n�t��^�Lc(�����#S�d����φ	n�ĀMo.;sDZi'<&<e Z�E9
�ũNcF��W��<u�����������o2����֔�i-�X�lY�}ٷt�N���8� ��O����֤|s`�`tP�q�IwSu<QM5=\5îZ�a����Ya�O�R��A$q{]�Q�-�Б�e�[̅-/��(�pk���j���{����O�^�ы鄄ח��m>����:�y(mm~�,w��W)o��^��NC���>ޱ�Iړ�t��ʯj���}"Ğ/@8�;ɍ���y����t?�yj��	e�?(�2l?�ʰf���^���)��r�x>� v�Φ�1ǹ�֨�vNJ���o�b`�H��}�������5��L�T��jOsr��B}�'�R)j�n�<�Z�'H��c��&�A79K�^��y��qO�X����/��NDz��"�=�H)���t�d`���5�j�f�j�f1d3�I��o2L<��y'�jD�Y���,��g�# g�K;܇��~�}6���M�+W��ؔ��W]Пl=SS�R�;R�H���=k�^������\i�D.�w���q�/�����3�%p�š"�54#��P�Q��Qc2l����Von`�>Fi�h5��=:[m��3ȩ�<[{b]�fKW��jo6h���jTe��|��x����Ln���+��_v�Á��+}�¢7�����8�ǞNN�_��4-��8���e�=�Î�]�~':4�Ϭ�W6D	nL������|��2�NSC��G� 6.AQ{;9�W���j���/B�����)�{2:	���xX�9�gkpI/�R]1�h��,v��w>�Et�B���oٳ`䓛C����M�~��;���^1��80��I��9�E^�Rc����
�ƹ�K=�C�0﷮�N�iuʈTG�x�/&�Q��F6�|GpOԫ�O���z% uQ]ʥ�����B0�-UV���gJC@	���-]\ܪY:���S
d�=�`i�$0�<]c=�����>5<��Zj�)��޽j��<�#�.x�t��?���þӲ��B7Xy�P��=��1z�L���t�{Ϗy���v���]A)��p� |�?;ܫv��Ɏ�ȮU�����TMQ��1�A=1*�.���Tf�U��:1�F���,�����|�=��y�u2R��ȕs��G(c�����9���l=^�u��lgI�UJ�b�T���0/.�&�5[Xӡ�7�y����33a8�^jj���P5�Ʉ�<ol��ĨV�]>�tz/|kl�*_��&���_y��Z,I�>i�L���}\�X�Fc����/�)6)��V��c��mn�9*�<VMn��o0�EzW��Ļ��� �b ���?΄7��y�!ݐ��}���p�+�K���-$��C���\��ǿ3 }�GW��o�e9�UX�s�*L�lF�&iA���O�A�	�ќ����;�l'��W��+}?8�D��.����rI,�J�E����K)�1����N�+s��ރ��Bq�tO�]++%7��;]%�dn.5ͻ%�Ԝ,g�6t����d�kt�)��ԯ� r��r$��Ne<.�SO�p���-^׀:Iz���Z�&��P\N(�,������):��še$��_��"�%ٚN7c�X�a�2S�}^ĭ�aO�uR'���x/����p�MG/�8��noW���d�=�w[?!���g�Ď�޶P]8�T!�=�U��k�R��4]	<�^�9L4�Y�K�yn�}�F�nRK��4V�,̃�S���]ݏ���K�I�QO��'TV�월�^y�0���q-JZ�e	0����,��\��.o�C���>Ș-���KJt&�E	���SS@-��OUX��,k2Hfҥ���6י�)Կ&ͺ\5L?����<�������t�|譭(��ָ1������2ҹݫ��У���B�UR��ֻ/����ɀQ$�3�^i��V6��!���8�|S�G�f�_��᜗wOg�V�7��4ng�����r��ʦڇ���Z'd[Ƨ�q!De�d㩿�k`�X�3t�$X��Z��� ���D�X�Y`k���s��'X�����.����h��rxR^��Ԥ*F����{��r��1$=U�����q��_�/�m����d�'�͏�bK�lg]z08��?��m�2��Y�
��N{���~����#����H�95����_��KH�pbBˮ����� �+�n��+-������2f <���ed�T��z��,+� ����M��^	�]S��	&�b��*+���g���6�7��S��[0������<�gn�>��ִم+���ģ�76,�ݎPi���*�K��3m$I�� ��~��pt���KO�?�AɃ�����8E���[I��br�X�ۧ�=��!�6����W��a�)��s��w;�p��m&\V��G�ľ�`e�~��|o��i��h����O����+���>��Gp���b���5}��Ȯ$+��ΉO�H�{%��;� �+l�JV���p}�W�H�2o���=\>8HG�K����Q:Q�`UM�:��s��+�2�t�Ò$��Y#��q�'��O-�Qt{��S��t���g������yʥ�6X���&O܍g+�zN��L��RfϮ8��׌Xz���bm" ��al�f܌�9����&�t����)�UXt����X�6΀YA����u�Vf���h1g�&�w+Qz���]�aLo<����[��gp��	S����\7(}�a���/�,�)
�e�gg���ǡ�-���E�mP�t���*��-N�l?�d��OS밖�D�\�[Y��2��Z��S�2�I�O0Uj<i�\[��������J�y�}ĕ�� �Ո��	��6g��2iY�� a'��.����ɥޔ���'r����h�����Xoʳ-�	�qh;8��߼�X�~�,����2Q?���V���-qRդמLI���؈���&��V�^��N;�����%��/�!j�Y��1� �)W�V�7"5��)�-u�[��.8�[��ȹW+���6e�?���)U�Q��u�E��*��Lּ�T�O#�d���<VoW�+͢�RB�c�Ďg�Y�������r�fF�v��>�.��_�`����p��r,sZ�h��b����$Xj}��$[d��"_+4��g*S��eƦ,^�3�\�| H������wM�����Go��

䧛ѧk��t����<�d��'��d��N��+?�h������w�ҏ��+e�oҗ���&���ČB٪�Y5����2���y[#JY��p��k�F������{y�f�a��s��Z����qK
�q6��N<\�^>Ͼ\~z@���x1H��e\|������Rz�g<]�EJ5k].��IW�*��g`b�\��.���ZU��b"�V����;v0��/��g@F2��?:i��	;������Q�3�d)k_���h� [����[;͈�-;�kK���7޲�D?���ݛ���K��II���j��lK�^&���z��;�7�7|;�yAI��e�"Pƥ��<�Ne���ۤ���5		@�`@���y�e��\s��&j* c9 �z���dO���.�) �>��M~�"�pR������d7V��=;Q
�N[W�e���T�8�����,�w~�_�4
��u�H��{����<��vrΪ�KH���b�ָc��Ƥs�C]Ώ�s�ϕ����1�D�{}j����̍՚w۸�ma��?p>��|��3=��I��t�N��es��HR��j'�aE2?�_������#�i:C�#�L$�j���vz�,�<$l�Kc-��u?�K�h��K�3UNW��	8>�U*JR\�!��`����
��}�S�ƭbÙ��BR���W�ӄ�'kȯlԽ�Zp\�ij�[�}�rc)��������T����09#mNیxw���iߘRE�֩�����̒%���gi�_�ެ�#6���-ϖ%���s��ԇ)��2q�䧸�EߗJk5�g�g{�N������A�~:�lʿdu�yEm�1 �j�Y�J�ӧ���=����?�Zg��Y�����������e20�����Y��M�.�E[��j�aC����.8��飦��B����N�I]IK�^f;���V|bwja/�xx��l�v	�#N�
l�(�%����b�&������ل
�����*�����/��8HA�wl�˓�kBR%�L�,�/��|�~�"K
����Y�,����|F��2蛡�̗ID�1��8���P#�x�l�Gޑ����0m&���|_�܆jpWd@���N��M�5u��w)6͊��,���^�L>>�%�pn����tx�AV*���r?6�M,�v=��/ٖdIߛ{XF��Ha/f�`w�N0��I�}l�Y����f�������gP|X\;݃��In���b��O��@�"�Z��U�ҵ�;_�DA�cU⮮}m	F�?n�MjM�|8�I�~um9q�?��q�X|����o>��=J�W�?7lI�i������m=k[2j"qe)�l�sQ��Sƕu�Q3�:>��k�.if�v���t����o<}G���J��n�r�:_����-���IvRE�(�G|Gz�����۫)oX��!�&#Í��[;
�<S�~���n�2�����IL��?��K�vs���tl+dkRjx�����Ǽ���$K�lb�'}@�K��n��99��'��T����~|�/֩m��c����xS�|�9C������Ѳ�1�G��iD�sٓt2����)W% ���U:�[O`��K�a�o�r��d'�gU�g�Җ5���`�
͐�+��D2��X��8K��v� �Q�tnt���D��X���#����I�=}8�P�*z��{8�R�RX0�̮;c~������e�tp�a$�����eݜ�����!˰v�:T{��H�\�9��~1�"k��49�����d@e��S���CfwW:	6��*(;�o��٥4kh��ˏ��#�����ĭ� �d� �׷1-��Dj�����f��kh;FX�A�O�~.��\�����������T�	$�m�$�Рbݷ=��&�S_ܯ�X�ry�C3Kٺ�q�3�-����MA�N���D|b�o�[s��[G���Zamk#; U�x�vֽ��&�ϖRlxg�2��j��m��>G���)�̈́�����BU�^�����'މ�����w�o*� .y����ј����[l�#�ֆ]�Q�QN���;4Q������P"�����Bc�
��!$�|�ə����kaI�vW��������/�������˙�ɜ�]~���C]	��j�!ppsy�s�5�fB<�MՇ���e�9�Ϻ�5>�����{+G��
0�>Ք"�h �ò�B�i�V��\�r�SpSt�ɺ蛱}i���W�P�Q��Q�S=K����o3SrD�</ي	�C��X��#�ѽ�����+��䩵����[�5��Smt��Zm,�^�t� �b�����jG��
�AҳZ�N!At�d�â��G	ؤ��iRP�im��[�]�w��L�O�;����E��h��|���G/�g�'��0=�����mHԇ�]>G�-t^K����r,�H����@C:>"g7����9�_�ٛd�{�4Ua�-y�D�Q$�;�9���%Pl�	X�v$��Z�ʧyۦڇ &���{��ZT���A݋ܿ�0�b��6����,Q�[-���[;Y��!�7᏿�Β[��p��-���JVx2�L�߅�L V�3(6/�5�{�����?{��@�55G��j�
�'y:;C��E/^*�d$�~1Ya�|�I��ĉ�A��?9 ��Y\���x*�����gn�ba�g���5�/�'��@�O�-�=�,�m�e�v뛹��d��D�ԟ*X�٫��Yk�>xd��h)i��#%��JA��:Y{��A��8�KAe��Z�6��2�597+)��J����d���ooo>oa>7[~AIII~!~!!^l	^wgs(��;�oܵv�t��a����3on���!{����J���F���J���\؊WP�ʜ��JX��JX�J\TPB�F����tz���
,����������#�'r�S�O������^��]l���s ^a^�G���O�[��t��+��æ�m�г��                                                �g��lX;[�rysA�~��'.��'V�O|���'�	I�HH����I�(/��Q�_��Lq����������������׻y�b?��	�)1)�����n��AOqA�.������y�+�FK�Wh�6�f��:Q��k��)��t���j�<�?����6���_����+�|�Y���z�ym�fH�&�)������GqŪ"��j@j�Ɩo� ����m~�h���[�� �[��*OL��v���c�j��5�9mL�#HR���O��3�Q-AI�ɮc�eC���,C�` ����3CyE#��7�˱b�uk�����-�N��5��D��U}T�u��H�1�/��1���T� @�21<
h��s�f�#��<8� �:t�n���8���1����>B��ӍF󴷠���<�1'��	������~�*?42���t}h9�Ƕ=i�m;��f8��l�^���#��w�5��y#=�(ʉ��@��x���h_T�X��:����9��:�����G�q*,'��P��_�Ȏ�:��c�qro�w��?�g3��ğ?1&������C�̍�Xl>֚�) ���6��fb��E�b6xc����f�O�2��1  r�GK���=A��f(&u�"��v ��]�1���YO|,����Z�{0@���)= �L��W`{�f��r�W"%��FE9������n$�+
��Xв�H���hC��0��c$�(Fc ����Y�A׌�MS�1p��YA�N-ŇТ��.�*	�i8*@V��qϟu�,�C![<�`�~�@z�"@�*��>l���W~0��u\������g1��ܙ
�ﴗO�W���Se�xh��9�ƒ<>5i��Ք����+\{��ƙ-e,���~r �!���]E��<h�"k��' Vhgx��|�WZ]ZZ:t_��G��/㺗!��	���5�t��B�4��1���s���
��hgv�Ldע�œm�-�;y`z<}��%�(�׬�PraǴUf�8q��"�Q�2X�1W��ܨ����\�c��Z�W�Ã��3�~@�+!�6�������+��Q:�E+2�JƟ,�+���%o�����k#�r\��0�������z���nnz��z<{�{�q��k<�O\���7�o���J��n�KB'��0���`���O�s�� )���7��kK;�g� <��i�P��t�MO?��c(s��ss��"�����q5�%�f��my�7b��N�b���ݣ@�c��"^�{|̕rdVf������o�\�%�� ����]S��Fm��3�b>NY>�A�\A�J���-
[P�jl[#
:X�炶l���2���(�[;��ȍd��<�ϟ@�y{���v0�l���R_ ��x5Z1 9��_��9��X��1��i���j�(Q|��o���F{���=ē��BP��EY=�������|��SFW9pn{�ǢL: ���*�\4�E
4��z��-�}�5����fjDq�@?C�B3#Խ�bz8�o��Ga,���������hcM�Q��w7�K�ڄԓ��|G�$ź�K���k�-�-�ܽ�;F��t,�5��	���6̣�mx�$tg���T+2*�ɝ��̣�,��I�奅�>���uz���i�%��g7�m��#b&3��S�4��=g��b=R�viO�Z��E��;X3`M��Lj'5���0[��$�@���O�>����*{�I����N�{���w}1c(�ܙ��(P�TMV�[P�uX�R�o���>~#��+���%:z�$#�\��8���v�j��xJن�ʶK7l��9�:�:>��L�L�����F�FZ-}9ҳ�&K�������Z��zje��`�������Y�1C*c�5="��:������f�L��E����
��Y��i�Ѷ�\{�84��#oݔ|D�����v1_����`�Ʃ_�^�ǉ��+�S��,�g77&�W[0 �����Z��V�Kz��Z�e0�ɾ�����.7��#���h��^� �0��fg0�%�U<[�}��~з$0|)�?ξ�k�8LP\�>!�BЭq�u�Q�>dZ!k�?g��*x�PT�e����Y��G���6��iQA;Xc���1� m̖_NYJ��5���s��Zm5m�H��6n���I�Wx��r����=���W�ˇ��E�	�3>e;���Uո%�B�u��B����[� {�%shڶ�f���#4ő��W��(9q�b�!9�O2��t�x�o���|rfJ9���AQr��-���a��ŧK��˴�L6������(�^ȡ�y�����Т�V/q7i��֋�U��� i�Ն�� �E�g��D�4h��"�˧��Z-Gl��3��Y�Ǧ<���g2��B��������7�#̮wZ��DugϤ��^�,�_�oo�Z�m��4��R����"-b�{����E­Z��Q��1�J32`�`Iv����$g8�b↙�=�f�N�tW�d���')��%P�{��S��\�M��3���w�=�}���I��.���.�{Sy�����_&����9<{�Ư�Dipg>���v|�.��]���fRu��"����6�����?50�` ]O�%�jx8�Y�ɧ���b��m��3i��0 '���+a��N�<'�g$^�R��Qa�gN2�L�S�츓��ĵ-�ī@�e��D����`�L[NEj���6�r�}j�d� ݲ���E��{���>�_��"� ��ψ�N}K�밺��<� �ݘ��1��x��_����Q�"	���%����E��4�ɕ.�m��q_^a��
R%
����M�-qm�i;<'�!��~��� @!�C��4�&{3Z�k�\���T4�h�b=z(�B��5Ub6��*�+]�� n0y!�Y��~��Q73[�T�`B嘈0X��)� �4E�$��Bo?�p2S`iY"��w&��;�9�&H[R3��-sA4��� wڹ�YW��$��TKw;����UV�������Qri�hΣ�=DK�+*��_�6�2X��&}F�avj"������m\9C�g�����!�O�M��d7N�R�e$Nw#E�]4G�d�����Q~���hyj������?��8���"NǿP:��
��t�v���^Ϯ��K�0�Z�K��M�v�O�dm�=�?�l����L~��-���r0�:������I%���[�觺˳��CVQhHlf��+doҬ����zO�I����hң8�w=�v�����?�\�̫�W���}�O6;]Uk!��6������]�=,�k~�[�nF�L1D�w�ꈒj("����?m��K�eKU�?�zJ�fh��O�4G�$�(�X�~S����V���>c�%�k�+���p�^u\�������ϳP�yk0JQb� m�z8��H����L
�O�?�>���V>��ϴ�ta�.�r��}s��󄕴��~��2W��}����:�Mf���X�O���u��،�~̐��*��q�/��^M�ɝ�bîC7�,�d�BºzG�p=Z���_��ܓ���)�p?�Id�1��Tv�3"��%�bH/�}�[�^t	1�M�t0l7���֭�ۤί�	Ԕ�7r �0���Is�2	����YW��?+ t�g�qEQs��H㲽�o��ף$���}U�rMfB�ӏT�=�.r��fF9&d['+|�뢾KQe4��fe��k���3+Z�pYz�L�%q�H+܀�.F� �`!(��u�o�%�O�� l����1	����]��_H1#_�U��1�*�i���Fh~
�ѳ�h��5^��܀��mg@!��ʃ��)[0�Te75j�z�iկƾ�ht��Խ�l1mt��4끴��F��Բ#�����0�[k�0��q�/r'�#i���w�Bf{�?�(�� ���r��/�I��1��`4e���i��ӓ���Te��f��CM�%�u�	hSÐ�I���%���Ӆ'(�����z�z�n���Z���,�B���<��kb�Di"2�mf��۱U��Ї��elu�6 �!�@���̎ȫ�Χ%J10KS��eЫ�x�X�P3o��!(nۃ9��]Ԃ���뽬c��\�=E��pȲ�<8#R� ��:��~W2^j^�b͗�P�-��G�H���l�n���z-zZ�3r���;�;������dY�����p8bdf�)� /|�`�q�h�
�f��aBҖ�譌Q�
cE�v�B0��~�<�G �v2��S�_Ļ�>��[��b�|�r#N� ���x�3��L����ݰ��!��˚�ȱ��;X��f�w�	0�u41�3a�en+Y.ɞ4$��v�0�þ��7pOFKR!�f/�l#r��7�������-����%OՒ����8זo$��|*�2;���7cI��\.Xr~ ��Z��J�%��H�94�nH.	����%ڽ_1����+U�6
"��d1=�j�:�r#DY�	:L�A�[��{W�}�d#��*�;R�ܻF�zXoWR����@�͟'-r��Sߧr�.��A�:�j���.9�4��Ew�ܡV���!��<�Z� 3��"��1@��Մ���kx������v��sWQ��HZd�	R!r�>�A��e`��-��H�(��o��Q{���枑�M��������6��tsW�;�>��b��Lß����`=/mb�7��?�'���j��J׊n�����2Iw�HF�P���b��6�ɞ�S(qCj�b����A�kf�e�����4�۟�Se����gyvy��9��$�����2���Ghk>َ��<X�g�������������"��6�/��e!~����@-O>3-�T�&F���,��q��.���RIk0N��6�*8"X��m�:�ad�s�ۀ�/1��NC�t����vR�-o
_=��?��_�	|�Ҽ��'�0	�R�������&�	�ׄ�˾�67�2�9����fE췳��g4�`&vu�9I�.� �C�S�~�+�.��!���_DjZ�#SS��_0�$���ʋf��o/�m�h
L�\����X6u����B�.@�Z��D3o�R��C�V�Дx�J<|�]V]icr�x���U���"3MM�����#��Ob�J��E#��-G�ø`XFBf����;FǬb�W��EzR��uY�UI^GzȂ���q�"�pZ�.��,��E��%��ֿ�,� �E�#�ᴚ���Ҋ@|�z�DhB�A&5^���	����&^��}Z�)�ݒt4\�ؕI�B2�]���t|�QI��p�9�*g�sn�꿚f=�$�����T�2�I�󟀦a���0��zAV�{��n��	�*ΰ&X��1���6��C&��*����f�gV�M}��?��-��Ί�n2ق߇#э�󴑇���ഡ��Kx��f�:����|t���Na:���u��I3��9�q�u���P��îv:��=A��Q#�nE��%K啶��Ȫ�$��`G��>�'�)72$�.��N=!!��/�t�V�_���0^L��8؋]҆���k2��V/Y���j�c;�Y�UL �Q�� ����f�Yd��xKI��=/����\�D�{�����jQ�jOl�.�1W�7�:/���ZOW��M����)�jU�v�	��c��X��.�=�?j���[� ��M<�Ɯ�����v�ݡ�!��I�N�����?�5؆fG�]�PF�(�|y��c>4��e덻b}OF��e�Ζ����t�
˓e}֣Υ��7�h<ɺZ9g�mi�!���.��Uv����r�kV'�ӝ(И���o"�k?B��!�B,mwug{tK���8o0ۄi��o[=�?�P����LԜ�(�o�/�1�P�[H���,X!��V.��m�3MC���	����q��q�秏����x�Z���O��p�O�6T��<�q�UJ{�[x� ���Ñ��!X�9,��'oymΊ{8�Ak�(>+T�|fR>��<���y-���*�l�U{�Vu�,��%�Z#���giݠeP�Ј���9!�a��t;�6SH@˦�C���e���h�Rg�������W!;�F��K������ke��%bх���ݠ���6�a[�n��B̍�`s\#�:<7�5��/�
k3��E�
͙�^)4�ॊ�WY�֛e���nJ�]�?'���]��E�&�X�A+���2��L,'��z�Cʪ�J��^+���#Y5��/f�v
Xj7��XҖv��D�]�:%�D����<��@�A	��8�JFx�\C�q�"Tu��}g�l�ʥ�5��W�s5f�4�7?~����b��i�@!�t�ۻ�CAr��(��v}�'(M���U9ڭ�1I��%�����/6M��3�,��am`����*A[��~�u����#�<��:ٖ'+�Fn�y�nC�L�*	4�M���5�=a��@�	c�
O�>��ܸ�M����K��%��5K�:Y2�p"׮i�o�"�/Z2je�}D�H�Xd>G|��_O�-�Þ����Oԋ�����p[�]�p�y5f&���=���l8�E�ck�����D,�t%^WS;TRi��x�<���ژ�f�8qyM�g��H$��Qu]h{��b͸sC�+iv�FE$qli������j+��Ӊcsf���Y�%�)���a�$�)eI�b�i��.v��&���PR�}�O'��a�#d������;��R������'��V��~�Am������zR�x�8Vb=� �#��'?����+��
Z/�k]��8�ڰȹ���]��Ƒ�ձ-~�wm��}c����C[�|;;W+*���>X�*�f�yַ�L;�g5��D�e�N�-��H���>q�H���E?&���OF�Q�;�`ffϐ���kS�r�wg�ȼ�z���㳛����dܸ�s�i8���Z�5^��M�6˧*�8:�D�%�<�?e�v\�C��4��۫R���V_6<�YP��T���s��x�\��{d�K�GjDt�
�T�{�U�DA�EΘ1��p�]j����G�m�=��ĩƺ�S�&�&Y�9v|o���!>����ꗌ>\8�c�#2��l�kg��~��2���3c=А����ۓ4F��H��RР�-4|��3��=���4��L|ch��x�i��H��|�.�i���s�Sp�ӧ��r��N̰����̞E�/�����������������!�V½��ɚc��|�l��5:ɳ�K�o/�r(�'v˚��=��D?�ޡ/K���Z�Ş���T��uQ9E��<q����Y%+.�ީ\|  
�s�ux��%�S'0@�m��q�.ms���&*���O�����Do��>�����g���߹����,R,�x�A�c���U����\?y��Y�ā�GҖo
�~���9n����o@�awl��1��ǩ�S�&�ic���ǟ>I�_��X��LCZgOo[��3��q`O�\^=��I������/B��6��	_�Nm��9G��L��sNˇ9BM��]�zK��u/�|�R��TX諴,���w<�^u�uD��p�v������iI?�G�#�y�]�Ǘy#��u�X�u r��4�B�;.-h�BxJ�M�+�vN{�Ī~�@g8�]��LbUI>�G�N�X����a�'�*C��|Z�	��R�qZ=2JnvM5a�y�=b�	
�Hb�M���I�F%a������,���Ѥ���ҍ�CU�ly;��%�@x��r�ؔoP�q�Ȍ�V�#b��q�?x�|/3;���I`�w ���}F:"�tQ@!�Ɗ�P�]�hX���^8d'Uw�ڵ��>K}WbQB���E�?�S��n�'�����kF�����f���r h�������3��!u;ڿWS=̯w�1���c l�K�ќ�KV��@�9ߌke�����&y��K�h�M>���<a��f1^]�8M�� !�嫯�(P�ؤ'v�z�M�k��v��l%�oN�F���U��7_��]c����@_��:�_�w�r�,��?$K�(�+������I5V\~<$�ԧ�V��%����*�ӎ��݆�y�H�NV;3*��C��vm�ʏ��ȥ8=]U��B��Ƀ�h���(�AyVFdb�Fԣ
8,�HK��{ϟ����m�`GG|��x;��*���z����ː���Y%����k6'��݆���pD�%������{Lp�y�Ob����o}��zPz�=K'�j��Ǻ���P��#��D�r���C҇z���;)�_(z\�(A�B��(�_ȏ�X�٣!����ށg�~'���p`�[�Nt{�"�����g�ϥ �o��u)[���T`���'����Ĵ|�^�|�����:�p}+#���`@���\ǈ�������<`cI��5��g�uj��ZlS�'�a�\����"ޗU�_7�W������q�aA���o˸.�8v�QG�{�e�qҌ�e�#��-���emID�-wB���C�J^�(�m��E�ON5VU	�;AC�q9ܕ0������N}����M��3�����2�qd��zmW��$����������S2��
��X�<+�nX����h��}�hK+����h&��S�G9_u߶��J�����B*۝5bF	E�}�"�b"�a���E�e"cd͞$kd3Sdf���~�����{��}������z���s�|��|>����:�k�\R^��J���c��� ��hL�H�5��g9j{�,r���^�Z�q3��8<�2����)��ԯ��?��m��!�񱀿��_�]���#���Z�/�i��4�gz��0���ύ�V]���T�5~�W+{0ҵ���V4� .n�ܓpF��'(挰��_�$��_���C��f:�vC�r�ֈ��q�%�l�VbL�%}t�z�@��~�o��[����{��fxk�NU2D%��,��u�����/���a��o{ݍQ�|�!�:��qsTc ���ʭU�*�tx�l'��ǎ���;g�.g��h��ß�_YJ��}�"��25��Ԡ�Rd{@��j#�U������IzRd����9��y���H��Q�(E`�9m�����:�M�����~]GRh(�������G�{��ve�e���']�*�8�ۄe�P���>�'T�Eݣ�_��,O{�)+3(���!u�l���`�I�R�,��&��
�͛�_�:p9QY �#�K�&5�j�	sp�~���S�G��V�~d�K.��P��H��#��Ζ�p����Uo�����l�j��r�l�mW��硟�F����,�>)��/��8�����`bB;M�!��
��Mrh�+�!�0=�P���v�{�O�$?W6A��U5��暤mu�����)����ԩ>A��}rt�ξۣ�m���F.T����ӓ3{}7��z|p���ђ�x�C��'���1{�b66Ę��lP;T�Z`�h:�$S�q�Ɲ�Nus�����n=~�b�@�%2�.09�T)�U2Z��;�	j
�k�7SS�L�eݤ^����PÄ�։P|֝�g4bђeNX�0:�+�.��)W��j���=+9XU�W��s�I�����#�V�p�����W#�4�%������w����i�>�mL�#�t���W�4�\�>Um���c ��f���A��)��x�JG6"�-Yl�	�N��ݹ�ۓ��mPF@�����-�H��B҃˦}h���Y�~0{[>�����n&;f�@��66k8��&O����|RO|���$���5��T��S-'����o5���Hӽ="��M�O7�H��אǲN�"�_��4(vNk:��rJlm���Ǘ��\��p0e���8�"���+S2��(M��˹���Z���ʤ�>�F�˩S�A��y7�(>r��q��C,������m���V�_X@o-㺐Uh0O5�3�祚s���h/C��c���0��)��t�YC�0�޿d�Y���	�&u��B<�m�8t�jH�P�?P�BQ+�������Ζ�#��>��Ż�)Vxg��s1��>ń.<����P��1�����D�P�����kRQ\�V�u�oiN+sȎE@�gv�[�lÈ��2���֬7�-$U�2�J�qٻ=���11��f��k����bs�G��+����S܏�h�=�܏4v���m?ښq6L�j���5~�0��rB�<�y�; �9��6�@練I�9�Q��~E�W��r,Zt�w�*��ܴ�Fӕ�+d'��|�.-�u>x���x�������F�
�@\�XE=�`�)Ї/A/Z1G$����;��ݭ��(�e�Q8���Ȍ���^���J�O��b��)ĵ��d�i*�U����QUq�)��)�`�`����#�о�R��](�<~���}� ��-�|�L�[�����O�Ѝ˂<��RE*�E]$I�pK�ߌ^�j���\��C�씐��L���{��r�6z6��;���X&(�e��慨W�շƪS����<}�&�{p���"�2�((�"��&��0bq�Q��?;d��:�)��F^�Q��~��I�ي���%�c�|6����{A;��������h�.t���S1]/K��<��(]w�T<**�f�UTmЦ���k8gl�X�6��G�JS�9�sI<��r�F�چ���'cp��{T�`;z����c�ig�z�J��Y�a��"��V�9���]2�ִ�b�d��9�8�5N ��4�>�o�#:]�3�Ғ�`j?_���� PGZ+��:D�P�ȯ�"�Ef��_<j.�n�dȆy�8���Z�ah�����v �)�]�3N�X�\�֧��aJ����=�`�ô�i�@�b�#��V�\�i�=�7Y�$�C�J+i�7�$��8s������T��mj~ 6���S��k;�i�w���x���Q�؇����mŖ*�i�B�󘍲̄��*?j֑{��o,�Nfl3ˢ�4y�4B:�IOdGۚ��0�Z��4(]�t[���o4;!|��ޏp��E���_UK9�=dc�nn+g�5�b������(� Q�qy�Ҿ���-��qI�����ǋO=o�%L�ƿ� �p9�I2�Ci%4��qH�b����<��Ogy��?~,+L�Wjut���P,�υj���^�w�`�NH�d@��(?l�=��^(%�B��t�7T�3$��y���,>����M���l���v�@tQjR�rH��IIq�;h��2�'���G����h�,�n7}��O�J�]}p��>��xb�H�Hf'H�CB򋣦��n>9���O�}�߼gxNx�2�W�fX�y5�?�OE)m�����N�R+^�~[�v�^Y�g��6�Ͻ���u^s>�q��jFj8gk
d��-�.t�{�n�o�9�}+�n�?��ݷi��^&��j�������O�X@�B+;:���q;�D���y��m�9,��Ef�MZbbT��9�x��*�X��g�{��#���遷�4��
�.�15 ��R�r��}�M^���p>��p�5rq�+�q�y�W�����=�m\�5�C�K� <��p�9`�=;l��PQ�Lj��O5jU2�꥙�.�E�� �@�Jbj�u�Ϯ��L+<�xyC���)SNj���SiMp؟̛���~�|)�2����\��9��j�6��*��t�S�͕
=����.�.��*B����5X@Z(E�g�~<�Q�"�6-�ټ%Z<F�	��#�����.Z�Q�,#�ģ�_��g�/S�K��/C���]��,��}f���b�����o#V(��G,�5Lؐ"�	��a��R��/B��H0l)�����;'ޭ<�;9z��J���������0oW�c<�Ԏ�����A���g��tti��oe ����[ ��as5Ps[!4�i�W:����;�Z6`�/�߯�׼6i6ފ2ɳ�j����fHoc��x;j�)L�I���-��G7\�ֿu��-ȹxJKu����<7})�휿hՐ�(^���;m�p��Gы�s#��a���$�')��dh�mt�b�N�o�f|"z����.+�u��:���I�ͼs���#��\�Z3�VK�oj(0���R���Z/��=n)1���u���G�uw��س	�_h���8L7�~6��㣞�雐ac$U�m�}!"�0��=
s*��~�Ɵ�g�]j@-j��~�͍/�]���,�5AE��"�Z
ؤ�DdW�#�*�?I�S�1\���$b#�l��*M��JYS��l�J�e��Rr_O���ۉ$G�q��b�!�D�wYBKE����"R��w$�GW	E����#��k��F����;�`t�IaF$��S�Ln��wT[�2��nTa��L�Ϟa5~���nگ-uh��w.� �^\�$����/�nXO�r����`�0O�[���e(jv�hB*Z�.p}�$`�%�u��N�?�C�P�E�bj�z��-�����5Rxtz&�7��7?ٓ��=���f�͠���j-��jV�{f�,j;��]�������}W?%�#�u�?�r�:R�'t�|8��0��<�ܩź��\R��7D7t/�v�X�?ie���u��\I>�F��s�����kȉ��ֻz���.��_�1�*2�q���bi3P-�~����mLl	lT����D��\�]H�^�������7�^�E�j�R�a�N�!N���g�V�'p:��݃8�(�\ ��B7�A܉w�fW<�xթ��j����X�z�G3���/���63rY��Ҟ��̾�e��PYe��iɦ�k~��mN�m̏V&��FS�TChW�B6Ƣ�:�S�������T
B��R�P�h�E%���|^�v���+��Y�I{��܊R��_#`�rSJl=�"�c�'a��]դu��7�Frq⽲Z����Y0��~_1��"����4��Z�6'Ո�3%#�(𸪊i-��cg���9[�XՑ�g�ߩ�,��Cc�ON�9ʐ��P�G���Б���vNa%I�C����x��=cD�=�ޓ��	���*�7,��d��E�	�A$�E�ǠR=��x_�g�$!x�����3�Ү�~�w�m�Ƭ��+��>�P/����������䏐��tF�drj��]U�q�B�����Ώ}F0�vT�����,����ִOq�X���@�kQ�CW���DNs*�?�������+6�t�k&�NU��/+���rп�eS��58��C�ʝ��ti�s9�-��u8����^_��� YCۭ��9?@��,����ks�KM�.���K�hf����2���ׅm93��]�fܜK¶�55��.��g�S��q/��� ��������;��g��6�f�v��]�$ױ��:��8,�+�¼yX����`A�����>��6�1���}�.��!Na�O�ݯ0�y�)��^jNY[rF"�
��uh�.1�����>l�6$Z��bg��ӈ�䱧���>5T�XNj��o��!9�	rݫ�`Q;BRؤ�;��U�׹/|��Ї��=�ƓYM�sņQx)�I�����xT�5R1��0�JO8��i8��"�׾�%���lT��>�����ż�M�36bb�`�f!���/��Z��̎�c���w���@U(�z�'}�i���3;k6�3�*S��`S���ǔ�veϓX���5h8۪��!:E�0��RL����2��AN�?��w�?�����2إΉ�
�������8<l|\��cE�O�c��h����2S�W�l���s<�7�;�#eY|�]��FY�ê���y,�uR���Ĉ��(��������T�w�#[h�&y�Qj��T�hy���Z"���,@�] ���3��U�����R�u�c�l���#���_�W����G�7������G�x��킩�=ԟ��] C3�_�F�-���C�;�#�O�x
ǭ��çħ��B�)=�����S�oS<�4Jn��*���K���Dս馥ͻ�z��lQ��?lYX�ʅg8�/,:��32˨�7krhw�16���V��W��S?�M�d
-0�ځD��n��x�]��!��Œ	ϣ`���#uʿ�1�v����լ+���t����<;���
�X���H�����Hכn�e�[Y<��S��TN�I� ��iRn4:����0dz7�a���W֮q�DtBr��%^ȝ�O�b�Ya9�G������^$5M���U����sh�#�>�lnW�.{�H�	.�v\J��ѳ�h���v�xo�"2q�w�������w��`A�>䱦����}e�"��3��~#�*�v��D� �ԋ�߸j>�Ĵ萯��ɅK�	ke&�0J�a�!a�L�����j}jy��1N�J��ϟs����L1?X���W�,���Mm�l�E�`�f�Z5�֩�&N����o]o�yO�#&�2������r��2�o� '�:C�v�?���^{,��v׳�=4_��ttM���s=���GW<�|�~wd�!`7���B�Bf�N����p{������!v��[+�8JR7�$g���~ �l��W�wP�p�665f�����������=Ǧ�)XQ+�R�����\rK���D�K��U����+3O�+�L�7�r��U�8T=�˕-csq0�gL�vp�-d���կ��_#�}����reTb�đ�a�t�^����/P�*����a�5�?hFCvT9�������H��R��4�F��Q��l��`/n�����F�˘�kT�K���;r����h��hYyf�Sc~�[S�����:,x?H�v�A�Xj:���Ӥ�jqw-f�L��;#��ᅸ��o�Է?��tx�	�b�UƠ�XpH-1F�'�>}m=m�|3 �y�$PQ���!��Kx������hUz��<?^@.����+�W��r��x�?]u���Xɝ,ܑ�ӁZ������Nz�4e>���H�%��G��}���>H��z��m>�����z�J�v;^ӸJ�=m�y5�G�ӎ�g@������W
�6Ĳ�1e�˵T|��Dψ��j�]Tj5�5�ȏUnMz'y9��6�FJ���X�<LW#�
�|�[6X���e}k����ȑp��_(~n~���9�)��琶/��ߎ+6�\C٠��6Z%�������5��!���C�,�[P� Dz�=o�����r����yo���;��jq~��_�f�\��������Ҳ��6SE��1�֎n��I�3옮1�s?��lBy�f�E"-��V����׭;��؋�
^)��} mdC��B۠����x��#���8[���МT�.d���F[3�VT�FP��%�Uex�� -ƕ0~����<W�R�K�F�xC���^a:5�i�Ԏs���,�q.��
2���*1��	)ݠ�ct;�U��3'̖�M�����N�w9� �L:�_9Q�k���<˭�o5t6cW��k�DFU(�p�]���WEұ�:�V4����"�oǏ��8ק�y��k-l	�-�l2Br���hJ��Y�Rİ��KR�\б��+\7�L�
umr��R��PB�mc0�l<O�Z;�y���sHG�[P��?�سQ���C&���N��$
z�� Or�/��,��cߑ4�\����WkL#���D�PMf4iVz�K�+�6�x�k~*���T33����戚���X2Jx�`my��E�X��x�v��I�z��_��P|�$0o|8�̣�r8!�Ϊ$��0�v[�jD�q !ɉ�h���A�~gѣ�gxA�"�!!B�**�� 7.h�w�{�t���Rug�r�R|�H�����<�GtDU9((�qX(!n+%A���pu�;ɥ��!�0�O��$+i�=�E���Y@��]o�ݑ+-�n�[����Ŏ�H���W��q�o��Y1T�x�>�ۀ�>Q����U��ʞ�	�Ǥst�Ӽˤ�{�0�Z�eWX y����-i'N�A�bR*��&��|0bO~�\wp��oܴt2��+��L�!5�0I�������6Ɇ7�*�Y �đa�hg#�:��9�$���F�Zb����;<��E����
����C�P�a�<2�`�8!�d��L�0u_�w�kːp[ع�#�rCv턂f�
`����jw��U�r;�t��A�=L�+{K�S�|�&9Д+��Y>�7�x-�2�=`v���4�yl��̊g<w�$���d��gx�m���V3GE@ɛ�7kk�J9� 杘ٵ����_�Q��GUUr���O�&�cg D���!�u#�=�����6
r6'g���jdC4i6�=E�0M,-�V<Y�Tk^���x0/�~���/=4�->����(Iٟ��/���ެ�)��������[�1f����r�y���A���x�Y�Uh5n6}�&3�M���#��O���ZY�o�L6,*d�bD�m*��_N�1��_-�j?Q�o5��{.>�&���[��j�X�M�1l�ys�� M���B���wM���.�z�
E���[/]�P�����$Z|���ݧ�7����P��#0D�H@tZ�8B�*Zo��\"�vV*m�|D�8��{s���!�W�hv���J�Js����!H��Ί���R@�\�W������y��b�ѥ��t]��,� /՘ȵ-K�		��g�"�3r��.-N9H����7>����(D�*�W:D4�仿��m6Z�Դ�ڶ`�n#������&_��k��m)�,o;��� oo���(� (�-K�x�P������o)MlPY a��{Nr��<��+�UU���NT����)�����#C4�δ!{��ߛz ;0��|^�G	J�j��!MȌ�8����A���QE����`n�����Ķn�g���3g����L�UCv���ɤo�1��{���vb���$�p�NC�V	��z�ߙ4y1����}�4 ���r�9y�s��y��/A%ؒ��)γI����,`lD~�O���g�Ɣ������qX��3�4��~��c�x)��cb�5\��(�BJ;+S����sJ$>D�$�d&��M!T�}�lh�h��i��#S��IS�@�����_4��FS�<�K ����S_�x-ɟѯm�y�$\8�|J���[��9���3l@���N�F�b���GTm*j��,�fg'�#�l���-��Ú���yqv��~fr���:%�?XD�_J�s uGW7��olVB�f��^��;�,}�C�\d��G��!�Fr���D�T׬E�1��� x�uC:����x���'x�����'��q�r쨏������[Г�vc�W�6�tK��O�̝�@_N5�x�Wt:Ɛ,QJ����%�/���|��J���㟉#��e��~v�,$��2&��(����jm�g��}B}Iq��7S���aA��"���OzCv�z�P�P�ݓԊI����
YP5p�-2�=��7��6��j��5[M�ЕG�x�U!�J��F.6cʟW��:u�q���2ۺj�_�Wn�����������>�nE/���2^W����}��Hg�I��н(J)ڷ)�v�5�����<���,�y���^	m�0�`��`�a��:9���\i�
+��퇶.,Ϩ�ڙK�:s�J���s}��\���� WJ�t����~�����@�B�?re�X ^��"��y�))����^�0Ri��7ϐ�-��c��S:T@XHa*,抍͓%�&�e�y廼��W�k�z��tܝ�{\�<�7��;ҠHkX2xL,L\YC�S�M]��I���7��&7�����;�#�R�[��wI�Q���	p���I��KC�.џ��
S�}C�N�H\��% �H�i=TDF�Gk_�c@ob��͵��Y��^	b2nY\ٛ鲄Æjg���	�$�%�妡�)����=5�{��$�J�{}r�o����'ȱa��pڙC��ʨ��;y�j^"����B��6���rS�2���,>N�\�B�F7�Ρ&[	=)p<]F��r(z���bQ��6]�E:��Br�֯'�E2�w��JÏA$�.*�Z\_t&�$���T}�Y��ʿ���P�n�ړ���k�"��'�����%��-�j�S֣'�GH���9ʾ�j�N��m����apͪ���f�졬Œ6i$v��0�5�{6f|+���h?ψ��9S��H~rwIQ/����g��Zֶ'�HǙx���On��Ŧ��%�>JpC)��f�"��,vD�RSٯ��[���,�\���F�{F��\����l�ꩭh��_�[�u�a���fZ�+'�B���	c]�5�q�����&��K�	C�p��;j4��:NE�����8���T�6�E��j:�_�c��3ɰ~]1l�+�Ƈ������fm!dZ���'�Z��&��}Z��Y�œ�2�71�͌����i	�JT׼x�R�9@7�9?�<�l��k'���E�!������,�\��[�&0?q�Ӌw_��w^�j�"�P_�:Z�p7ac���E�%M�S���D��췱<��y���H�.�r����䗠�e�^'��}{��<AUi�F�Kj1�'�1�����|�ԥ�{TM�g"�ԗ��E((CAؾa�6���Ӑ����#Ҍj/��m]L���7��MF/��a��u�J{0 ��"��a�t�ҁ�(��ݭ��xݰ�F�|Q"r��q><��7��K/7��u�� �藨_��]�����hF�ێ��6�`Vwt�)	k�	��DGc�C)ӡa>��);�fSSdp4�Z�#�P����$H_���tN6�M���8KO��g�q��X�'�D��`ǣ;lF�7&�X����r��ŋvtN�mQ7/� i�;�zOd��: �\��e$/wX��6�c1�Y�4���5g0�t}D��(-�-7 ߋh�W��AF� ��Q�Bf��(H��>m��[a>Fu�ҽ�(��f��:��\�gᥨZ��0��@m-��h�:x�J5ud�u)�ۨ��i2�)(�JG�q2�5�8�FH!�v���E��׀� 	�چ	��7o�s<��������4H�u͘�D]0m͒�������	�:�,ݮ*l����Av|7��⪪Y@�� W�w� �O� 5����b��7�U{S���h
t��p>����j������h|�q���ks�����_�.��K�9�^�{Ư�5� PK   �beTT�a�f�  ً  /   images/f9879790-346d-4fb7-a00c-c72301b216f4.png4�UT[�����kp
���.
��kq+��[ܵh����	��Cqw��7cd����>k������AM�  �()�j�l� $E �������EQ�  ���iٚ�  �d���r�t��<8M��I��^�k)P�� �\����}(�R��(�E�/ M��D"}��[���P��X+r��4�x�	ǯ�2ٖ;_��U���*���7L�W����hO�LՁI`TF��O+�c΁���;��pr��\;fВ�p-�W>���ͫEdp��{���err���t ��k��!!�?��1��&�����D���FƓ�Ҿ^���  %��a#�љ'1P�;��sw ��P� ��N�?�͎U��@E�, L���\|�fe!P.�.����377G�p����;�N�|���� FL+�ZQ\�`T"���|��	�`��V��I��I<��+'"�u�4M� W����B9H�2 ~����2K"����m簥��U�pm������v�9*I���)����Q�x��'��>Z���_��)$ �4R,p��]����Bb�[nz��-�d�q���k\�7���7tqO,��u����ZR��{�g@
�Hp9��" �3� \~��T{ Ռ�%��U�#ts�K�i�MM��Fx`y�	�� I ���t'60��ֱ���nR�T��U-��d�q���7����׵�:��v�_|������(�{o�G,�Ѵ��̩��΢��[�3��3�z�$FN�<3�e�����t:,;�	����#5F�gȺ�)��ǵEwH<Ie����
n0@bn2��\�+�8W���0u�B]�$]M��-��m�����
H��rS��>\_~n�xZ5��i�%Qׯ-��ׂ7<浰���##��꾷Mbxii�5q����~��G?-���a%��Ȣ"׽��.ISx��Oj���=S'��?>K�gf��P #�a��A�R@3�c�����\:�QVF����Z��.��pn�}(�n�[��ȉ?[�_�*���ן�Ԙm57;�q�C[���~A�~�h	X�8��yгW�j�P�0-�9����������;cy����>>�عd'6欽눈�wy׏\RZ
>1J/���q�)Xf� �P-es�����?f��7Pџ�,g�y��555��"�j�SO���ߙ����_̹� ��7�~Â�'(��][�z"�a���/�,�x:/5�5�n0�YSk��7�)C�1Q�|Uo�+����渟���~�ڕ�7`��!�RH��#KN�����Wx�7=ǁ���_NV��u4�wR

��哥p7��Zwx����V����F|�����=�����&'+�v9 �*U>���/�{zz���!V�����3r�7{�g�7��]�ihz!-�1eZ����x4O�:��V3�F�
����a��_�ۜ�"x�l���0 /��ĥ��7irۺ9�X�Ex>��=��Ȭ��|���sk�a�Nq37����(�&�^�ޏ
xd^��Ѭ|���;j����\�6X��N�WX|���x~�VWS���G�l\��~W#6o��w�kH�O�R���b
q��;��Og��ڮ��sWn��[�rJ�t����|.?S����2^:����)�9�����'�9^n�^	|�.�����#�
}�D�.<�E�����y��Qq�/ih�i��a�4%Uy����>���� ��v���F��ǵ�~���9�b]�p������3ƾ��Jgw��&���K�7б���cv�ԃ������,;Xii�����hv�����s��?6�ۡ<	������~�Ω9-H'oϛ_�Y�A�.�hV�����hi^@�!�����rq�4����F�Y�go#�/oqNX�gZ�c�{&�A����~;"�C(�)ʌ08	�w�%S��Ƶm��̈R걷������'�ȱ��7��ؕ	��%�$D�1�Gu(%e.�ՙussVl`�l�1nZ����RP�=|��iۙ��]k�H�s�z��طz�.��޶[۽���#������1�#�������ݵ� ����8ˊ �4/y�;�=�F'�ۭ���"�	�ˆ&��i(�~��X/�������g�狮�%�n�"��H_ ��@^>�y�G����㮼C���B��Wuf���~�б�y�:��N7�/�������]�{��R'��b'=/�؈h����8�B`p���Ӎ�p��H��_�U٣��:�����(�t��}2���^t\h�nYs�~B]N�5��Ͱ��y4���7䓵�1�{B9���2Y-���qI�c=�L?�_[֋
�R�>~�h�|7�G#�w�(T��d�8�%D��E��#�Q>9�ŗK��"8={�-���>���oݜ5JtYYYI�/=?������ل'�e���f̸������������� ����JR����䅦���˂���&�[���6_�'N{���ۦnJ@���y�W�=�H�3<�ma��)g��T"��x�3�I�΃��O:*�B��B���!��6^~ �TO}�8[�5��)�c6���(����k)���EJ�����qW.�Ğ�=�U��ݽ�^�9����)n�c������l�3b�$cK�v�	�����&s�bo�n����V���w9�V��HՇ���E�f(�)�̧�V
���΄�dR�����g�=9cU�9�)N��}L轸�Q~�'�[eƻx�;��s��h�i}-�����oje\�
�������YR��3j��Å��߿�R�dfu�5���F��7�揣��P�K��?�+�٦6>Z�����J��RNO�[{R�"�|i�IH�5����		��D�� �GT_���f�˥`�I�&�&�&�r󱾜SZa��Z��#"������؈��ʙ�UmIII�������r�#�M��N~p�����x�L�-��bi�Pq���B�/�����=l2���b��=u?۹I<�\�&j������������l����
�ɧ͘#�Ŋ�>�O�Q��;�Y��`\Qۅ����3#E������րjJ���zW��	{�{��Î�ߖ�]Eъ�K�y,+�/F�.~kY:��B�<q*��� �;�b����K��|�v�-��C7}{	P�A6�p�c��ߣ~'��KAA�K/�r��`�z4��7�����]U��S�����?������{gG�:�p������Hh��EL^U�r_ѨL�V����ZO�?��ǎ/>#n։�~L7Bk�<�I���????��������i��ؖ�}Ւ��o"�,<<^Gw,�f7�EO��3v|��us�z��C�?f�K�����q4�/�C�iC�J�x�=}x�j
?дsa����Fx����޵{�]����eg�%���0j&�KԴ��YI|#41�XG�X�1ǧ���v�9���svu}�ijȁ��ݟJ����˪�q����,�G��Y�ex����<�M�K���_�^�� r�7f����S����F<�,���í�a"-��/9���v�rQˆ�������ʙ}u�˿2xb���Ԩ�&� 9��λ��;�k�i}���X���m7�;���og�@��jԻ��ԁk����%�Ep�E<�������}����1��x�#��K?|CK�%�@|�[#$B.�*)2�����Z��ǅ��wO�/p~y�9�����B�׉��Ma����_z���}�������m�֛��t-�������
Ot�϶��i[2�a㠝�@�rxT��K�n��:nGw��^���~�n-���ԫ���7K),�{�|��{ˎb�����LJI��2��JNv��j0��*����^Z�l^	ی���|fk�p;汑����íZL�E/��n�冋�c�����u�����EoVC��}����a�W83F�� �
��mĺ�Ԍ����(;��������mMw�
.�JWhǵo��ߏ���<�M��.x��R2��5�������<�݊���nGl^<�W�Ŵ��(a������^������SQ#M�YAO����!~�h�x_$��^;-�Zm��.4:Wi�`t}m�m?�~۵8N)ej*����g|<���X��;�ﹹ�-n�)'O}��d'ǥǆ.r~�Teע??�_u�щ-՜1����� g�|���yp��#> �s:�%�)	}��<^��@Bc܊��=�Z���J**�c7�(��A��E:�Gq�u�j��a,L�vg�������A	S�G�h�,%~��3����=�'K�@
@��A��X��d��L@����(��k��ˮ�a.q��Tk���ki[Ī�Ba� i��:�4�d"E�V�Jb�V�bMͧis\$@B0>(h��6��`�&�~���ж�'Eh3�Lx��oȒ��P�X��r9�Cs ��D)�Q���Zʣ�"��wtj;�ɲn"��+ذ�Ё��� 0*��A�{�dH׼��n�S��!�.8eg�Ԕ �a{�-�N]�o�C
Yp0�lVhGH ]m ��d�t����t2��
�h�i������D�b	�tn�|YfX���&v�W3�����p�p<]������k~+�]?ힲ)�p�!#��I�X���j: d	Y�Y�tEEsyVhex1s�H&S���gp���G�.s�5�ܣ-),Z�Y|�❢�uX�P�a����v���A��]|�t?C	(�@���B��(�4�}ކ/[R���?�p����4�;����>��p�t���m����8���O( C��2�10C �Z������:�W�BT�(�Z��?�4�Z������q�S������)�Lw���r�]"�H�}X_!����v���qݍ=e��K�Q�F���X��DO�"s|�6VĈn.��������b�U��ۓ�e�y����iA��_k�����k�HS$�:枋t��'��9&�PB �!�;�Y���8GfA2�肼g����3����G�ǁ�?�RN�=׸uz+��Ȋ�k��4	�L�g9w3�yF�TД�8,��l����ݹXS�@��LZf`Ep�ZZ�|>�6!��N�ʣ<]b.�h����y����.�I��	׀���*u��J끔i9�.�B�аZ�T�~t9�8A"���A�n�����dD$2D����絹���A��(�n���@@�1I����6;/����������;*G�OX�"���B�1�֫ܖ̨���\Ah�9�}^$-?%��Ϋ��9���f��w�q�!ʂ'�qm�>[eqr�		}qݏ�M^�wx�	�?SX��I�Ĳd0��i��3/`���.#��#�-b�ш'�1��<mh77�d��hu,u6ҌU�1��H����|�c�������>x	��,;��� 8]j��c���|K�����F�<�� �EY
��F>�8.�%�T��Մ���I�;�^�n��6z$Eg��C�H[;���:k뫥T�}T\��%YEv��ҳs!H��J�-5���_].���	��1��V�`�A(]��h*�G�{�U��޳ �>M����[��W��@�	�oM'��d	[�=�'r�Q��:Cg����Q�w�[�:R+JX��*�C���mз��D�Zz�U'7����<����ρw��O���B�=~�~�ki~`����9�����F_�쬽EV^� ��_�UĊZ_��\�B����Y��y�
D���W-M���@�!��(Q�Y\҄J���{�L��y"{�WXMb?��	���]�}��;�v+��4[�+޲I�h��cB��B�4;;��C�c锌��zU ��3���X8�©�[��S|�N��{B���Mϣ����1��o��G���O�8�suJ���\XKhH�\, �n~��׫?��$�z�����
)�f�_R� u��2����"[�c�g;<%Yx���;��: m ?@7�A;��5��x}�n�+a�o�a��>I�R֗f�D��}F�=Tu��ʜ�����}4�w������1��I�4���MW�����[I�|�O�M�"�^cܴ� 2��ࡩe*�6��)6
 ��q��m�V=�Ŝ��٥`����L����'Rz�Ͽn���<�֎���`h��$�x W.�`�ST��A�.ګ� q� @�;5b�k�4Ukg*pYS���?9��ǭ�����ɚ�u�@Ѡ�4�� �$�9X��Vݔk`���S}K������a�H�*u�E���+�Zl֒�oF���ϖ���l~,��U�-$��ۏ���*i�q��H�hz�rl��N���.:V1���&[|om:�_�O}Z_ﰚشCt����Kb���jY��`g�g�vV2Ia���~�lWN�E��4c�v��eǬ�E�xE^�ݣ��@��ruJM���y�#����R1��� ���T%�ƈ�F��l���.o��g (5����$F[��{#"�qb����E���.��A��*�.�fA���$������Ⱥ͸�|ZF��k\&�H��V���T��>�-��u�s>sr�s|�=�
ֹ9��NY8�/d�e�A������,�<Q�ta�A�LU�W������W|V��o�cQ#���B�(�A_�'��u3�ti���(⯏%͊f����p*��˿���>��������ys�u`dA�� �C������A(�x;�7��β6eHp�$Y�B�,�?�\*\<\}��'��o$
,�N����,�l*��);1{^��uL�;���|��2��0�{{�'��C�eP�#J|��
k�"��Wm��d��_����� Ƨ�L�a#��ӧV�{���ڜ;P��e��w�6����{9f�9�u��hE��C~��枿�@Tž��[�2�6�-uyYiYT��_�}�����������p��"�����m�:�Ӽ�ޣy�.=nk�����ZI��	"�>u�܏U���%_����XG+�S~�=M��cxK�7�)����˲�:%�� ��u���9C9<\��C�ذ7X������6�d[�?�7���jڿP����by�o�� �X�4\������D!�-}����H�yx�=):��b��2T�`��l������Q��5�7�=�7�����(�}�
�m�������.�R�m��qX]=��(odV��iO��ug$��0$��C-R����1�9��o���sK��?(	}�sbhT@����9�.��I! c
�Q�n���0�.��!���n�bw��������I͐T���ǲz�U�.+�8M�`�7�2(��+�Rd>Gp�mb�r�݊=���ƚ	8Ri�������e5�,M�B�B�z󒡠�� ����I�89���S>2�v�� ��  "�����6ٱ4H1¨����f TVI�l��i��%�!���� {�$���G��}Z��lσB����)qKt+b�T��"R��m�� %U�k����cF�~K�j�j�L3n,R^����1�yK�ăD���|���h��:�cj��O#��د��$��CP���R��Y��H��b��H9���4�
iU"-�F;S�oz\H̝+�ӐHe� A��~�T��5���_�Tt7g�ps豒�	��vf�31�$�16_�Q�p�:B�i�my�߅w|��P_�%
�ɬE���M܋_�]�Rt�;Վ��1��P�IP�o
c����u�b��u�@�3�8���0�rEi�`�{\1(����5���g ~�ӭ��l�`��un@�d�=G(!����u�%f�n��#�"Ap��A_�&�ǂ�@Ň/�"FZC�1�?��M؈D�R�2[�f0v�����B�6iw���d^.��a�������h<�M�!�7�H*�q��'X"
��;DR~\�!�+�oF"�$����ޡ�)�����i�t	�Ty��P��5GXI���9��9�CP�:I�O�2� �
����p)�E7񽵣d�崳X��Lm ��dK��J��.�Z��/�ƶ ����m��������ͻ�Is���c�MU�pR�@���)@�bT��<���˛_��Zgƹ�r?xj1uxw��ǐ� ��1%�hj}X�O5i@�V�*���� �k�?�Cɬ���,�H��n�S3�抎i�r�a5FE"K��_N�N}r)rk���Z3�e|� �f^�-x�ɚ�PX�$����vwcuw��P-Oh&�	k��yrSյ3&��2��I�Bn���$�����6�׫(�DoBu�C9 �l��U�e"�Rqn����:J�D����fץ���jd�h�-�}d��S�I�UU)�-Ȣ^"l�M�2�OgX��x��#���a#�)ߪ�%2�i�]q��c�9���z�����w�-��!�q�LSc~k{�{8%'Mc�W!5��C�J �H��'<����i�����Ń���^g��@~��Z��}�36)�LNCc�=))���t9�F����S��ʲ�7�`�c1H���R
[Z����s\j�N{�a���(]CH�q�J����i�$�H����,%k:���� Փb[;�]n5�]7/\��200Z��� |�zȳ��4�:�=� H|@�% L�A�H��',bLv���}���yN�M�Y=T�p(��ɤ�i��\�0$Z��Xm�g�Q/�x���"������u-�4�d�t5���|��i)���D+�L�EZ��(�x��t�+N���:�i���Ü2�\@�?&�;k� ����bC?o��i?�h�Zx7f$p�b�3��5�j.++;\hԙO�Vd��O����6ns@pI�����^��}�'v�DM�q��t�(gMK�#=ش���OP-�p�܃E����!0\��4
\�!���b`L�y�F���OM%L9�$�/1*��[��� ��H�`ծ/]F��q����7
JYv�H`ld����_�_����lr*��x�B���X�2J e\K�us�vh[?�'�}1�S�9���f���V�g��"gw�6cy����D�@*L��?�fu���)���!�	�N�N��z6o��.�Қ����l�+��i2��ʨ�?�*�˧�X�u��o�[�!I�����N�p��6�c�Y�TxH޽E���0`E�(ۻ-���]"<�xj�K,둋��&���ɐ0�0���'W�t��ij>���zwa�Uw� �W���ؙ ��"���K�c�Z�^G����n��FU����p���1i�����@�����z�����R9�f� �O�5X���#���F��V���E`��וS���j�+�d6m��r��&]$��[�Iv�2�θ\׆�/iI�r���a}<��-���ù���v��:;��mG׍�+�6�6���(Ol�5�#ȑ��~ui"5���7֌��q^�L�XS3����ōYӹ�,+�%æfå���#c���.=W�.cg��w�WZ���%
�����Â�ʄ� ��b��}�+��qc�sl;%y1y��
�d�A�]�8L���7=҄|J��A�u*φP�ȔHF} ��a�;�f)������z�|���[vzO����-�5g^:��YD%���*�T���@һ��-�ų����*�����f���Vb��N1J6��:����M�4'+Mcrc��Vzݶ	�7}X�>.�t�gz�#&��`�~p��RVaUe�N�ǣ���Q�p�!
�=�`B�rPq��G�
�tf�K͗�q��Y�v����x��r��=J��a�g����)S�D)���0�?��!��A
l��K�UR_HBP�&+�Cb5Y��������j3�t� �I����f�����ƌ�6z���.�"q�NG���'��H��?�6�4�,�#S��K�
�
��B~�
��Y�%��ʨ�XU�����|'���N6 Nc"�D��QᾺ�B�����kOc���8�?���Q钔�毑� #>+qC6��W˺9��b��Te�v�h�>�vY�9f4��F��Q(hS�������0p�f���B@}�
jB�,d��V�2)��j(˹9�,v��_�?=U�Э�����=Tfu>���0Z�H?�̽�7RsP��&O.�њ�5�� �+�!�K1���Z��W�^u{å�昨�����@.�H/gӉ4.qfg7�%s��ǣKM�ŉC	K�
ӂ��ӌ�����B�8eE&�ϝq�A��I"�fv��PE�f&�|e��)�h)d�0�ݒL��?5���,f�V�L�'�����S�����Q�i��tyl����!�ƋQ�6:3��?�ʂ�^�7�֋�PЂI?��A�Ãt�fl�12��A�(H��ͨ&%#�����\(����,���Hw�P	W��	���:C\�;d��x��U���}��~,��]��ܝ�1�^0 5�l[6,*��Z�t�p�}�-}!�{N����N}���w�8�@(��+voo7�-�Ӳ���P	m5��� 8�?!M&�1k����~�8��K���T�����>m8�t���0���W~#e�,ɸ
�M�@.읉hX��d��g����%�~�*�McqY�����6���%,U:E�ʔ3�I�;���O撫n�S�A�z$z�����bd{�JW'v��[�Ngq�6^,&ksb �7�Ќ@q��[�T5X��A���c�6,�2{]�"�Nؙ�ֲp��rj���6�1��b�lp�E�X�|s��ڄ��jw��$WAFc��R �Z��DI놴�� W���@EpaY�����1cB[K�E�m�t�u�s�O��;����v^�~Sn�z�4$[UU���{9�p������aXK�� M��~�ɷ�$������n���̞maąy�[Q���s9��Ⱥ�n�oQ���R#<�9���2����}#����y�Isce:Bj��KQm9�"ُ��=K%d�)���P��П���Ҧ����G�������?�F�B���\�<J�e��$��,�vr�5��r��첑���R�-G:r�8l(��������찈�K��!���SfӟΣ�QAQA[߿��D-Fu�;���/�e�?��n7�2�����r��U5iQ�X�@`�d���h��i�d۟]H˴�N�Lx�+����jO�����=d�0�b���0��0�hΑ�%0�T�ۆ�M��A���F'2e5���!��#��DX�z�Ҳg��l��(!��dàb���:%����6)���׮�њ���D�V�_3����F�M����!�6�=P262��O�CI�i��0��(ͯ���$�5֦�c�8��_׵_��o�N}�*a�BA����� Cx���v� ��+w�R&���g��"�C�r�}��6�!� E�.xÐ���hZ,æ�O��v��F���_�	��3��t��$%��,铷�+@�y=!�DY�yJ�z�����r�*��2݃B¾��r�J&��Ǘ*�,������b��Y���?�T�f�m�@��6�U82	IDݞ.o5��Efy!P�ld�Wf�4q�G��Sp�r6�F5�U��k�7|�e�^3��t
F���et�{�^)T�#�$@lT�<�b4�nf�T�]Uo�� �`�'�z��b�=��ߖ��Zl�psB_�|��Ţ��lat� �B�>2@�$bW�g����}1*lia����f���ֻ�.�d9������'�Acj� ���@�Z��lOh'e�SY���a�e|����rh$�_EI��S��O��ϋ�� �}�rN3�h����"	A���<����Ho���XU ?љ�3Q2vH?���s��ci��%H1��� ѷt�L~�O�?3�B�ܒ��SQ����Ox�K��0{\||zB����W��Goo��C`��� �Ê�7�ð>m9��]5yܨϫk�v��=�#ַ(�����\�Q��{���i��,p�����r�N����ׇ�@���?	S,�u��ٝ��o\��d�D�o-<�|��\��9u,r����W�&�ػnh}�� ��n�����"���0�&:=���Y�& ��a�9�Q��c�1�+��Ӹ#j' El�5���h�_�qA�v9RG�$���wG�rϲ�c�7��;m��rt<�Sv�گ~*Q^��|F��E��i;�����< �m�r�Zh�-n� �q��%Ib�֪���xs�\\�,�4~'a��[,�;խ��p�8���H�6����j�h�����(�<�6���o��?��� :Zzd���|��A%ּ⊺
u9�0����s#q��o#Y�Mkwu�����x��1T��u�"�/�ʆP�fρefj�/wE��rE�`Z��'���㥰���G�Ix褹܈�[�69�N9+�j1�+�aT��X �T�G�O��n�&�(EE���x��~H�~�ta��;��pRs�*����eMΨ�RR�MS�`��Y0j(�tڽ͑�]_����,egį.�qŤ��(3D��BeL��z��$j�t�уH*�'�����h���Ra1|���q���	B�!r��Z��,���\�N��~����L�-
|r��D/hW&����\~+��#�_�!��o�=̺͐�(9�9S#�r@Y7\^���M:�P>U4�J����d @�:b����y �߰��Iy��[s*s^j�5�W�,��m(~ -��������y�Ը�		l�S-~��+h�YYO�����߳|�j6G���n���KI�;�0}�8���\v���˟_��'?)�2ˀ��̗4k}�`y_;�;��"���;��n^�ش����P��i��FAd�O�&L�������'��!�\�o�m����rۼ�/"b�Y�"pe�I�<�����r_�fq���D��j��Ddf�Kva�g�>TS�F�R��e�c���'w���i�A���w��R��.]�JlF*�B�U=����N��
�!	h��β�]gX�e�e5{z,T8���>���N���w���t�����K���cv�S�I �P�������������Q��x>�D���>^�!z{�AAA\����n��=Ɍ��������׊�T���Nw9Zjq~~z�()�����jy{�3q�7��9�<��77��˼��S<qq��Sm"��M�V-�o�gy[l��h�-��v�R�$N�<Wl�rٰ,,,�7�}��K���h���j��{��R8�L��˞]z�_ۨ���˯E@2�,ί��L����bg$v{^�Ԡ{q�ݺ�ǃ���ir|�����Ҷqr�X��Ms��+����-���OU#c�G�	���%�����k���z��V���Q�*�|Bi%ڰ5 mJ���Z���v�����1B������} �C�PG9���V(����`A��Ur�r��u����"gSAݬ�ӟH[�����)[��￴�XةP*�_3��n����� ��ps�P��5]������<�>��|���}�j,_?�@i\��c�/����z���w緇�-��aj��"R<\�ˁ+�׋��p}��C���ʟ7���$`ŏ�*��`�e�[��!p�{�P2�����^t~��2�^�h�H�`�𧖽п��/�́{�������i�`f���e����7�@7��5<��_5*�8)�����LdB�7��!�}�_'�-?b��Y���%҄b�f�	M]ZqU��8�5R�/�^�A%^��l��@\+��
�S�YiG�\��<2�����O�E)��^x�����Q����s�ǳ��%�e�ڮ�>�)6����M�����O���n_���2��ߝF��ʹloL���Zw����H~}�rX�{�!�!�i���������g�l$O���؂�`��}f�J=��!L�ʼ,����{���8�P�>�l.ޒ���jM�jvBjÿ�p��x:-�����mī爸�%��55�}�ݼQ�1j�b���m�sdd�X6e���;]>}o�\fo�؟f����?��̆��I�͔�JCn�V��a�	�F�C�o)Q���s[����ش�t�|+�@�A�0̈́|���`**��%�\�ny���׹	���f���Ɔ-��I;:��엫��3&Bg����ſ��;�ug�,"�}.3ݏ[�^.>y �aY��C�F�tz9c\>mG��쿛�xV�0tD�R�TBG��z���,�)W����@�k�1�g����6_j��D1�����!�!*S?�\�us��7c;x4�K�%oy��9��������8;~k|��:;X�����.�y~n����Ӛy/҈ �C!����`N�8 >��a���`����m�L{e�6����|mk}s�7�9��m�3�2y^�#�7��=n�lм�G0�����$���g�`����^ri����$+�@Y�g=�y+���iOٿp��h�C8T�@@B�Ľ@G��Aа�6�+��g5TI��J��a��_F"��!���OW����ʨ���}/��ݡ�����w}�$�cc���K�ގ;Ӈ��fn_+'�J��(bd�n����XZ,��#���;���� ��g^�\��ĭ
��_V�~�`��%�}�l���������(ފ�����{4�Z�#}[�z ���D�a���R�����Dj������8���-z��w��sB�w�#}s8��I�)�Ӛl{�zv@�	�:-��_}��Ь<Q�u�6c�˷���U~���!�z�8*�8�д��]y\�"Ir�cJ�u8��J�`�����4�l�Ѧ��'B>�K�5�|��֐NQ�����u��tuw��V��?p�V40yF���g��A�>F�f?=�J���El�=�X+�ϧr�J�<��T��<�Ғ�F�%a!�`�WQ�h���l���y��e	Y*��L�C\ \����k�:�@��Pt��J�ս����������?x~׳��M�5Խ����4��[4�K+LJ���ȴ�k�����<u��iY�s��b�̘y�`�P0k*�7U�j�d���VQ����I;�zA�����39-,I�5�0Ä����5ȕ�Q��yԺnr�5��Ԥ��g�*�!�1^�`�l��L����7�-����%�����2����{�T�م��</�Ԣ�KByu|�^���;��K�%I�D�o�`' ���������	q��i;��i����I�)�ӌJ������l&��!��߰����e��
02-qZ���oH��l:�p����R5�1FU�p�Φ}�a���F�գ2�*��%T�5o�ʥ����O�X۴���3�m�-9配�R*"i
J�~	#�Bnh��a�1hP�ˬ���#;T�]Tn|����O��9`�6���M ���@��v{��1Z�L��_�Z>g�#{d.]���\�6.��������$���s!�QW�{j����q8Ui��	XiS>������~�υNw�N�{�#;�4�LS�8�,�		�虘TjG�i4���f�q=,toZl}|�F&�2�xH��Z����b)�7(���%��7�y����<=������t}ؙprIzRY�Wh����cmK�~�����߼�$G+ Tz�X�	]I*b�#囖����	�,�P��>P��kπ��i�)�s���5sN}�Jo^}��r�K_V�%�S��,�X����Xwo"	��]�R��5��wf�
�;��Js"�f�����c�T�j���;XohZ�U\�u\\��W~���Xi���4��>�=�n�w�r��"�PB���Z�OM���j��'��@@������z��Yߪ�K��?7���ϫ��55��7���w[�:N�)�bep���n�
�Y�S P�/r2��&��j�s�ё�bqL�5�Q8�*����V��$�R��^�D�����`m��^X�$A�8y�:�M�r�`<o�>Kw2(kJ�tm�c��0�	�)�D��E`�R��l��66��<M����5���/*{�A(�J��.�9�7�W�]�?&��w:Ɏ��gٳ⾥�EˮB�?w�h��}�9�y��zb�/I՜���/Q��\� �(H�c.[U3M�b<u[���6�>��s��`�wO� �����n}U�Ͽ��p������V�s����R���"��p'�q��.)a�����H&d���*�c2ЋTg*ie��lI^Jp�!G�f�S���J���1j-��?]ߨ
�F�-�mc��N솣�����6τO���[i:�s���j	�!�҃�u�z���n��"�{3-�xn�\�7����7��� ��j���A	,@b8�Ee�v8mf�m���F����Bw��Y��5�qӱ�ĵ��mΘ��4G��\W��H{˸&��_|�Hi�Q�n�����[��DFOz��"�����HI�xn~��yp��~������ܟ�z�6vU���Ǩ|r4��J�3"�ϗG�&��c�~���?ʹLv�g$��L�)�%(h�U]����DVN�Ng��QO�QO�'Fr��J%Q9+b���a�]e����-q�vUlE	��y9��T�%;�,�&h�`�g�fʯ�*����Y��-en�6	�n�u�U�����<Y>U��SU��*e�0O7]���}�4E�nsf�@�@�J��M�������̙��v|�)�,����b������!�+�T��
�w&ݪ��Ekr��r|!ƘN2��չ�Y�B�Sl�ǿ3�zZ�R)!K|?V���ʒiO@߼!t�>m��4XxQ�r�iX�Ҿ��V�3���%N<�k2����2_;C7ƴ<��7��=3̎����H�/�jߝx������5M��YD�Nw�(���&g7��q& x��:ki#J"�f$/
N-|�W�/�����؎�3(�esc�(RFѴQ-�j�Q_bO�ѧ�_^|���^��W%��2�Z��y�|,�}��m�{b�R��"7/�لӘ��-��Xrr�� ���[9���s��a�2>ou�@MJ�Ӎ�R�ɗdQҰ�A�H�@��
�G�̜���A���<�0���<���k�us�������Ccb�W�a���vxxو��~���ر�/�?/��w4�gg.�Dk���$�ejmm\�h�N���R���8F2�|�"����JWQ|s|k�XO�I~96�M 6�[�9�9���PY5�=&�4QH�R2\ȓ�w/\�b�D��kќ��1{�}w� ����^.+������l%ou�d�_��B(d�@�A�-�74\�spN%�^��Kl4:n����8�TU���65����'�'.�~�6q~��:��KrEB�Gs��I���d�k��e���p��mX�F`�^n�v(�Q�J$;���qZ�5��V:̞ਏ�>G�̉��,�疲�M�f|🮟�XF"�/�o�s������}5�}��k_}��eBj�ݫ񍍍��� ��]�r*Ϗ]���N\�)�0�B�1m0w�H{��ѡ�a�ЎoA��\�=/�.��N*��D�b�����8�қL��~F9�P�������TW�p/�΄�]��&-ם�%7ŉ��6�x�HY�>��6��[H��Р��W�����#o����U	�J��ʃ�����|��	�>e�ά��-�E��䅮G��-0���V|�}!AW?T=:����>����"�GX�+��A���ߕŞ� A�5�����6�f�;�Hh�(c}0K���ΌX�p~���D`í�7�� �TJ5���B��Z�~��e�F׌ߋ}g�G�{�����z*�����ص1�|���w��rm����)D����!.�����ql��9pe��.��K@��a��f���<��-���bn[��7��o���:^N5���+S�le�D�eM��/�t��3Π��z'>��279���=ꈰ���x���}�6[q���0��z\杒z���5��/|R���6]w��Ux�S?�^����b(:�U)_d�C��r���۫Z2]@�#�+p��I��*������H=��)�-b5Nq����%kZ�}�i$�5�t�\��f��ut�o@I��Q �`��q��3�:��Kbvh��8����4?�;T��J,ij}����y����|�/�fD�X�&h��^���)s4��]��\	��H9+��SPh�.oNxj?�s&l�m�?���g4#<Q	�5?3
3�R� )�,J\M�YK����W&_w�h�Y��G}�ğ�<���QI��4����X��	xo��D)����l��|Ŷɬ�M��)P�	�hP��Z�>N�9N�9)j���4w^\±$�ÚIH���ĬnR����c�~�j�o�Gc��bC�顤y���tR:_�����3��ߛR��$m��9�Tl�?���lS�f�לּ��4 R̥�\v�#pL�sAj�D�~�����a�>э-GaU�X����g[�F	�2w���)h$���1K��1�{J��GO��"`�Mq���&;1��hu�=��"ēQ(��O��ݾ���:
��$K����e;<�vrˬ�k�p�H|�Q;�]jS�%���p���$/e�teϠd��Y)inZ�b�
q}��0�E����j��h�d(��p8��:Ql>b�s��k�TZ���qx��X�i�K�{͌:4�	��{�8��K�Î�rx&�lvE�`P�}�*���]����:n�2L8���2���{��i�YG%[�>�}�#����å\���F
�ĜaWSz(�qv	4fF�ų@����)�j�Q�0
L\P��
���|hw5NT�)+XO�Lo�Rz�?N�Q7�\!N��à����U�d*�T?v���!���Ƿ5UKU�U L��$��4�N�ý'5��k����#���(�g�`{�	=�W S���[�j�~�EhF6!m�ޚ�\
zI/��]~9'�st��o��#^��4�x�$fF���+�DR���"�Ԗ�#����4aբ��y�9���{r�bb9=�(�6T�0$�@��A�G��6�L��K�q���<�`����S1�.L΄;U��]�i(��GMh����N��O`\��t�J��X"C�(x�� -;�HQ�D��F!�^6�)�\��K)� ƞ�Mk� ^�,��xa
�l�B�G�
�Ӗ��%��sq�1ϲ�e���чM�1A�D�âa�1A`[��U������M�#�u�R3��R���ݳ��T��|�=X��yM/�n����ߊ����H��?6�bL�;C��W��hZ��¼��Au����9�a��r`{M��`�h�z {1��)�?�#����ՠm�u�������!���0�����ҳ��쨘�.��;v�+1���L��J�F�Iz��;{F"���R߬�EUp�۸�p~�!}������g�1��i�D�x�}X�E_�l���$t'/���m�e���W��:�7�Py.�h-���w�D��L��b��{���xKC�M����\����@t뢆�}kh"��pz�Z�bLo����JP��K@5�`��%"�3��l*ޜd���hgs������g���p��T��W���~����QZYW�u9����7��wy�(�V&J O�&���k����g���f/X�E#��_c�#��W�!���,���?��?�m#�c�c���{�D�;lSZS��vG��0�$��?o���C(�^��q��Y��Th�rX�	���!b��4dp�;��	e
&��>S�=��	��wN���%�P��v�5mL��N���HU
z3�W8�Eۚaؒk��:�F�J��Leߧ����jSgͶ5m�������rK��-��\�@��J,��0)AYFw�����"z6��
;����a���:'"�
���1y�	rhd�9�Pt�\�gͨc��{L�1ZV������b���8�J��V��c�Ti�� �_�Tb��tUGN��yRE�}|��dP�_�0�U�g�B�Ħ�n1���"f�̮")%I0�Є_@B��K�/���� �o�Y�z��`�؋l�\q��_���)�?҆�MTCU@,���$��
�gD^���2�ܥn���~F��y6钬��M>K��}]g�	���٣LI�ޒc�5Lrr繌�"}���"Z=��$T�[���I�̕���d3X�D�`�`,�5٘u� ��I�r�"$�ܦ7xWyǽ��^8�VW����~sD~��:ǋ�<�ɢ�#��]*�J�Ǽ�4C5y~>�%"��Q�w���rS���ܾ-ޭvuA���~?A=�v�Q~:p��y�)�,*�yIt(�����m/�ǧ�A'������[�������G$v�~
r��-;��t��~�Ԍ��[��L�K�8QR�^/����blܗ-��z��l�s����կ>(J�	��I",���J������ҧ��u��0��M��R���z�H�����?�1d#Z
[u�?hʰ¾rf|��-d��wN�}B�e���m"�E�|n.\���N�]��z:{<za�zs#�:��N$>@����'m}+I	b��ㄊ�������`�X�l�+�T]�s?���,��[�@߼)���}{��	��^o��W��ʾU��&�!����I��x�KQ5����<��;�8	�z���V��Vì��0�3�hH���&�EI|���nW���1I^:���ђ�}!�NST'	�PHIjȥ-�у}\���&������ !������Ù/��t���ˠvcۣ�ɬ޷&[�U�ΠW��a�v����XN5�"s]�lV�s��S�W�^e4�+ʪ��jp����ޝ�xm���u6��`�?����\�Y���G=:�)#N�;*Dq3�C��^aӎ8��\����Fse2i�!�K	T�T��Sx_ ?-�E΢q�H�@`��SH����
�?ӏ��\�#�KE��\�)��a,��mcI�%t�4؛��c�oX�i�h��6�Ti��1��r��w`6&8�	�[\��{������"Խ9`��is���cTR�0���I^r���t���v�SE{]Π�һ@f^CO%�]�J=avv��3�֊��Vl��x�W%�=d���Zd%��_��_�Ôx�Ǥ�$m;'olH���z�e9Ҟ���;ibF��
��t���[�>�ph�E���3��q�����k�oT-��.Tz-��.?���mӖ�u�x�/~w�D.yt3x��T
�L�Q�(��e��gY��e��)��
1�A
����Ï�DH�9]��+k����6�*�Rp�m�բ���v\h��d�⧘O�6�AK�^J�6>��_�w-N�R�7�¯(�1*Y�sj7�^�6�LN&�og��jS�zM>�������@BlJ�C	eE��1����\ąr>���`�YT>�pq����s��g�t���ɚZ�~Ѧ֡po���MB�7�\8��#�"kygv6,X��I���1�Ʉs�P��K�zh)�)'����H?�mx��&�l~����/_�jɵN���}�ϟ�rR��W��^�-w�T����\�DZ�y#��(	�%ډQ��@�P�B��0J��0�%�ә/R%0�aOfZ����*��`�j�,��g��.e�;��ZB�*��m)��h$�/wq�ҵ��S��8���L�i���	�����Îz� �G\�3GEL�l;�d�S0 ���)_�sIa������gA�
d�6ܜ�Y���:�}��i��*�E��B�i�n��b.q��4'u�Y�	�ĐH9��hy�����,ANj�pR���U�q	~��.(���Js��������"��F�l��WL#���Z�E>W��j١��n2�
X-5:`�j0���� ��I�6
U�"�,�̧��*�zJ �D�4%�?��E9�#g���9��_�2� +�ԛ���&@+�uy�Q�6�dl�x�/�{E�9��W�n��hKIl'�p���t�$�k��k�:� ��V`��sI��أ"8�/��d]"��j¸Ǩhs�G�r.�`�F=P�n�@:Y����z)����&7gF����6E'��a#�ӫ��P[�m8Wu��i�Q��J4ggѫQrSNy�j G0�?�V�?��D	T�A�����þ����3n��&=|�n7M�UO�"���N�>F�z5�`�5p�e����''\Ph�h�(���F�M�9}N*[��Ol�0JwOv%�=�lXC:Tt��KgE���Y�]%�Z�`[_�@%�2�,�s�[O�h�*�F	K@BR����{k2f�/<�⎚z;��ZQ�>l��rr���6)`K}��g5����pL��=�V��S N��7t�g���#�/����xR�R~�5�m�t�_W�FIʬ��|��D����p�8)��Y+N���k�[4���p��pc
N���:o��t���]�ߺA�;��d��4��8'�����xo��G��xe�c*�N��o��dy�ʙL�E:kW��b��:'�v2���ɧx�)5lhQR�'c�����z�O\�c�\6b��N #Z6\ߚ�*�LuܲI�w�����47�S��c��dZ]i���i��:�uK�U��&Gj���/��4�~I�����o��]�c5�����XF�N�:�q6˳�И�.7{�"��X܋Z�4x��Q�)�a�M<j&���)�t����X�>�!�"+��a�"xD���4��s�q6+�Y \Hg����5]��ϴ�_F�p� ����G�w�y½4,�e�󤎂�{H�K#��	�Xg�;4�������,.*�$�K�Tb�}��ϴ�BF�n;`��� �j�/='�����X*�~�d�����g��(ʆB���SJ:��".�\��
�})�"���5�}�ޥ{�I\H�f���=�jffH������9cc�+���ՈW�)�������V�p�%J	�*W@��#���wn8�sJ�P��5��#Aj�d?}�(H����WH�K���V�O�L9<�	.���W˯�Ua&����^v�/1Q��M��1�I\��-<,�N��X?-���k��#�q�3� ��C`\�8�<+#_��.Ս)?Ě� ��m�M�	�e1b��!'�2g�p�-�� �yܐZ8Fa�nY���%��f��
R��ێ#|&�������f7Z�<G:hX�5����U�y�~l�֘�<<5O;?��W�#�c���"Xُ���#�FJ��'�Q	.La�?8�A����G��%|.�oeo�D�U�����\�Xa��/�W
G�v�Yk�I���f#�9[^�?���X�N�ZZ��Ƽc��� ���ǽ�tr�c�)L�����&�)��0XP<�O�=��v��LM_$y��/��t�^���)T�,��9�Bn����k���rq*�/�6�ttt ��͟�	K�+�~���ּ}VðK���)-'���t�k:_O	�,fԫݥ�1���a6���k��i���f�D��
����G2y3��&M]7o��:o�3H�%w��gjj�����I�[�'�]�,lA���q���>�)��e;z����W��=T��#�eG�fO�:7�<�.]����:�Z����O����wpp��f�s\b�N(Io���ׯ_<n�Se��tB��,PR�]�BVD-��v+�"���ǿǞ��5b�A�$^�C��{��1�e;��a�ǟ�����(�_�ý�|r*�����_m��՝�à-R!Ǯ��r�:��F:0
���~U����4:�ŽgO��Vk�^��Q�d�j4�$���!c��cj��a%�r@g�]��t��l�F�գ'B�TX!ԁFћ�y�KP�������9�ϾP�P���'�j$OVǌI|G	��BY�����5���KX]���k�����㻎��!���t41�����EV��.��KC�4v��[�j����3���٭�)?���&����Y6_�o������ ��o��Eu�.�`|�u65�����;]����۫�>������i�����"����20O��Ҥ�?K��������&#]��"�)�F�	QoE�A�U�� �&2���2_��.�|����! c�͚yQ�;ޙ��e{����ijvN[��=*�d�+���6�Un����h�N�.$��7��˗�5c�ƙ�_�_��^'�T�4��t!��,�Ƒ��+J�HC��1uE!ܖ��;�a,���A�_�&g3�i]a�1�VC. �A�p�6EN0�x;���<1��eX�P�ؤr	��;��ƴ���7��	�j9�ٜ>�G�8Q"D����G$g�=��mɟ��Dν�n<�*�	c
E���'N��s4��8�����WcHϘ���[��]]��yJ��f,0��)u���u��}6)y��W�b�4�� �P��-?��d��ł@ү_�l�����7!��� �,�.L���Mk�mF�O��Q�� ���UU���yT8C����QpCCÇ_Ʀŀ�8Q߃wGm#�ia���V���Z����f�^Y����P�&)K����%g?�Ǐ���������r�	A 9-�Y�t"��,��5N!����ψߪ1�۫����}`��G�e�)�؈�_�\��GѧQ�#e�ڬ�1ǯC�]�����z�k��%a M3Q�IP���#A��YYy���1 5��z�\�S0��?#cFf�=�v+���կ���	ޑ�/����3�}��V��sA�y�NCֽ����s�m59�iUXҲ�����^��O�tii�'���VJ�3�_�����_���\ܶx��Rq�/W�Puc�W�p�V����n�H�A����#�[[��vR�>=�-���㴇D|�bV���m���!n;@�+��:�͍�߿l���<����E
�F�0���ԇ]~��n[��0������- ����V��3=?O��2��M��<4��� �v,U�u�8��
�xc�E�F0��Û՝�6�BQ�ݗ��ÿ���� "7���~)�
@u����.Zijl�C�Wj��I'ޘ��_io��J��&�x�˜��	�BCe߰�(�W�R})�H���A�?PM��������i�E�x���1A+�Ia�~����bW�<��G��ƿ�^i��H���y��^I�9����S�UM�/|�K.���ro���IrheM�۽����֔r��ffc�$��������苁�'ϟ?����P�CI�ӷ��Ԝ.t�ς�=V��-��NS w(&�ģ��7综ٯ�X���B�̛y�}�����s�-�s5J�
��8�֞�Ϟ��}=��⢠�c�d����s	*�W�`�����}���0w��������g_�k�E�2T\��悘II6��ZG�~7^|%�5b�y���F�EP��[y=FޤN�\�Q����L�P?�"څc�zc�f����3���V�߿i���k;�lhqozčfDУ9%�?!�6^����(:�n;��F�C��/9Qe����E���e��$E�s˜M^R�ш�N=�+r� ���F+l��B����"M��gJ��nؤb��p�)�~��W?�~�f�`����`�^:�4M�¦|!{��ii�; |"t���>�&� 11���Rs��?�q�d���fp<������t�Ƨ������b�r��K�ܶ\��FJ���J��b|��d�5��ne��఑WW|H��F�m�R��49(�4e���[�f���y�P4��j�,��s��T"Ν@O�|�U�zP�I,E2o���v2��c"c��n��YO�:w�{�{��ڴWS�r����^M=N��߿��ɓm�O�R2%�����M���Bt9�MW���kO6ߟs�eI�L;���0)	�#]]c�9�.7'�3�uaFḆxE�NT23X�|,q������xW�:꼯"�M�����Ē&@��,!��'h;��C4�� S�!?����#��I��G�mށ!G%V}W��QF�J'_�m�d�NO�y�� �JV�-��s�5P�(��/7~g�_i�S��!#����q��t�;�?IT�7�ԡ��x�+D$͹�ξF��Z�ķ�Pq������e����g5�&���ִ9���=�N[��돕6�0�����RގW�u6�7��$g�]}����7R�a�S!5�9A0R�N��?-����+���e�oy�� �;�:��x�Go;k�s����"2�c|��}�hB��_�x%�����OVMKi�ɲ���
8cٱ��Ǿ���'�q<�J`A-�+�
%�`���?���&�T��nAy�@l�S��(]�(5O_Q���n!�9"U���۬�X06 rűim���G+`$�Y��Kh����O��1��i�|���ך�b�al�2G�:�@,o}j��SY�~ʦ�6s�Gg���'�����cN0D<#����f7U��B��D#Lb[�����!�<<x�&/D�D���C���1�
���И]Ŏ@�w���@��\�4F�ym���0�eܰB�G5A�&��0��6(���\�&�;^qtR}�T
�;�:8#Q�31.�7����b�)'J�$�}�q�|�㬌2ZC���/�Q�a��1������Fe8�6S<</	����5R�}.�Ee��_H�^������������ -�&�� �:͑N�����r�1u���K�}zm��4��dK#�#?6��W�<�k��x��+�pK�͠��+Q.�.P���������؄��e`_j��#����*�2ٌ0��R��
Ә�e��8^�}1;;+"*�̒Fp��\9۵6d'0_���U[�~����]]r���|Y�9��ډt��]��� T�l��Vb��T�.Qn�Z��=�z4gݥ- �_�z�Q��N�}6����f߻�x:h�ç��7�H����`����X�&k`����:����_-Py�=Zl��(2N3.���C-=��F^oLt�ˑ�]�Ֆ�szQ'Go���U������26�p��lxC>l�_Tt�nNl�i�x!�S����"����	N��8�H)D����jb2#�����?�]�<�D��^)��C����ñ�ޞ$Zb�K� -�QL�!)�C��bK�۟�{��\�����[��&�o��X�h��8d?%053��I�:��u*����T~���J41^ �J�>��ܙ��?�u��T&^��D�����!$��x����v�Kd�q�Y�����g-[�vΙ,�u��ϯ��= ���$�������2�ElB�-�Y�Ä�(�a ������~����oSqqQUU%���T1�:h�)���DO/�ǎ#���	]�����)`�Y�Ԭ�6��������$|p?pQR� �b
;���"x^I5g4�+<�2�� ��S3��~^cmkkka� G�)��g5�N�ɗ�Fٛ O�7>�W��\Vsd��<�?���L��&!�M��w�WM�}�v�c��)ڛ'8������;�e�	�N%c[���)�	FpR�;cR����Z
����+PUX�b�����+Ȍ`M޶�1���"}$N�G�H7N���{��F����f�դ9�ɖ@l���;��LM�}��O,�E���m���ҙ������'
����zc��Y�`Fp8.�s���^�#�Ą��*�T9%���?29T0�kf8f�{�] M��S&6����涜i_���o,��/��}4��IL�Ͱ&�r4s�����c�2T�ڽFL�\�H�'lB�x˻C�y��`��1�YH���ߥ���Y�q�X��B���9�V[
��d��}�җ+����0f:6Hw�jt�<��f3��Ο� �i�%ǒ����}@��@3��@�D���w�\�R�$u��Jܪ��+,�4�Z��1��̼SV[�o�`5��8��<1�7��h��J^��Ǝ�����ivSM
�=�_TN�^�%�<�W�XUS�o��׾xXJ~�EN|x~yZ�����ղv�̐ݟ�-�M�:"�6X����� N�4����M{�9q*�=�M������+O�0��Y�P_y2�8� ��f
�x��jP����{tf&���t�q^���w�M��u�+x]�Y����:��o�r�_T��MNzn���`������B��X�t_q��[ZKa���9/�z���<�����鬎(\k���>LC�W1ɒ�-��ntI �w�Ja�C�NBBb�ȉ���Zn<�}{����Xv��Z}}}���tS��y��y�b�т� >	YH*����a|HG��jS��v�L�����k�W�"t?�%�q�Y�������B-��>X��Q����р���o��'S,����yfi$?h�Z|�8�����Q�#=G:袏�����/߃CBBdo�Re�6�F�D"sw��+	�8��:�+T���(���^�$Mb?�Wۃ����m���du�� �|���.�����$DD��_�ɏ��?)�^�R�}p�
�����S`�QY�
/j_~������D`���֮���gfN���w^m%~��!22 �D�]7��2P�⫋kt�%�Fs��:����������)����6��m��9`�ߠ(Y���ױLo�<�]xXXX\���<-���!zkc�B� �FFY���L�'����OUI�~ы{n�8����Hwa��ٝ�����+�D`}W�,q��/"~wt�Ƹ-7K����niiI�g�Ǵ�i �1��W2�{�X��{v�h7�I���,�4o=I����$��T���ld���#z�0kf�'Љ��M���{ld8O�9�1I�9{92_c��woz"x7?���X=��rjlm}�p�=��twL1Z�d7�6�Q�L̓�����������O,CC�t��/Wo'��w���|ֶ����d�-C������[�5���vn�y3W�_�q�zt]���������@WW���mq���q=+<[�`ugJm�8s>��ќ���`켿�ךit�]r�u��8:8��r�
p�(R�se%�B�����(��"K����i��ۻ @��O�к��Zᰭ�"E���>ZAAAr�T��'�΅ߔ���GCpA?�Zj����3���
p����͉��������ܜ�.����L�J,ݭ��i�#��f�W���q\�y Y���/�T�\���W+-'_����ݩ22/�E�o��b��g.d??d����>Yv��6U�LLL�����Xz�����$	����>[���*ljj��9��iQ
�ȴ��=��h>hkk��B{�>��;��l5w��S��t����o�Њ߂�L�֓X���7#DrԻ,˷�@�&''t饹6R�k�����W���f�;���>>>����&_V_/����01f,���Q��<Zh�;Ј_�z%4���o�+��eo��q� ������᡺ԏ����`Z;lZxy��(�x�� 5����W�������8R��ϔ*S�q7^�fYI	��,a�93^�\�0����Y��cmǛ��k�2�Ǵ�?:C��l���VV���W(���(0�cy��!5mmo�O���Iu��֞x�� ,���f���`�DDx^�_EӼ�b0�0�۫���{�%���>|������0Ofn��ȉ�����8q��:#�\UW�ˠ�ˠё����_&����
�yf��5otI�//������r�yȍ�X��i���+H��5GS;O����ˮ���{�f�1���l�L~+S���h^l�&pl���w�,�� :���z,G�d���ǽ�:/�=�9�Y����o;�)m;8��!�'|u�z=�� �,���;'�6���<�e@��� P�3����2���"�=�fT�h�2��9� ����ߩL�~;��� rt|*�T��� �"�H��|� MI	��s߾)�$<Rgzf�8�-���+�s�P���sk�:qS*�477(�3��V�x�pyO���.f>��<�s]��(8P��6�}�1�-,���E
���u�.t4�Y*�@� qn�\bP�|(Cͼ���%�P�����'�4�'WC�O�u
:^-
ifxZ\V����
���&�奥5���:zE��"�e�~ǿ�[ٻ͇q�L��f�����\ ��G��KM�@�d=T1谵�۷Q͜����ٸ|���-�b�?}����yyiy�k[ �ɼf��)���_����~q�
�}���m����i�;Cϼ�)�Ek���R���Xޟ��P�]X�)�	���, b�x���P���M$ �0o�:;Έ���I 2���L`[����9C���)U ���A!���3K������Qe��oO FN�v��m"��i�U_����|�����_`��[�O��G���y������ߥ���������Z)�H�`f鈖���ȎwK*m� ���ej_y��TVV��z ���;R6���V�~[�Z����-ʀ%|�O�S��۠���^0`�gg'''�� ��`P.�C;�y��s��{�i�HDg{3��?IG)��ժ�� R��	U }< ��#��@	���k��G���'R��K���I���d0
9�$���^J]����\	DX��03{aˀ��𤋮I�U7�o�!�w�Z��;�#��ېپ�u�N�D/��eT,S���#H�p~e%g� ��p, Yee@(��e���M&C��)���/��A�m�H)��ū��Z�����t��Q�t��a=B9� ��$J,���
�Q�=i4��|6U��t���!�0Qq�xк�~�������GL2�g����>��F����uIЏ�^���s��L���I��~�0�<��0R�����y�wij�����G�;������B|��i����O�j�x�`� �Ӈ�$?��� &�R�eKS+Nz�7��H���K;�oya���@������TWW���S�@��&(h����#d�o5��H�@�o��|q�N �Eb�c0)�Ŧ�r�咷�J��q��+ꊋ�K�-ҹ���gH��V"?��7�4Uv�J*zG���+U�oM; P����Ç� Ӆ2�9Nw��v�W��i;@i���L���E����ys�0��<���^�����4�|A�}"��|<����Ƕ��������0�@g7�|�;�1;k�F'����
��{���ǚVE�� n{��VZSCR�<X��r���8�����W��k���?��u�t;C�����,_:(�*�,>`(�`S������Ӱ4(]_G�������o���<q�#V�v�|� B7f',z���:��1�`����h��q@(@mOu�����������|˫0�	��G� �/ ��d�hL�EO4�!>�٤!4��~�C^�ځe�h��f/��?�Җ�5m��kĽ���o����_t����c���;���9\�UC#�ᕀ�www��ǵ.�ۓ �!ؗ���i�S��ѐ��~D�g~�0}��c�R���# v�������-����rmq	tJ[7�Uꆣ�9�s&�9��-r�0�!7g��:ZYm ��OI�0`ì	t*��=�w��6"�@�7�n�����.��}�������=7{B. kl�S ��&�F�/�ֻ=/�(�%��S��N�By�8?VUM�*L���*6��G�ۿ7�U+ƒ�4���c������M���+�� Wf�ft! ���Pڌ�N���+���G,Ϣ#Xb���N>p����} ��������GK7ggy�xĩ�����@-���gL�a�1���'��+ ������ߝ����|{���Tg~nn��'��-���5�h��<O�,��ksڠ�A�++s m�5���`���3`',������O�<</�$��B�����fEW�ۛ=Oq9p��~v���$�|����y ���^�@�t��O�cX���=�'A-��1���v�+t8����]>8�$=��^l����޷�G�k����=�j5	�0m���d�a�\��η!@ptuu �RC��$��r4 ���E[���Cl��.�&���*��)�} N �@?L�����!L��,�U��<��󀐵[��ٿ3������@F��:�w��)�7� ���=|�4snvV�{_�f�����,M���H�������00V�5-�R2����x��(��,����k �WUUY��{z�,tfi����~��V����,g V�#�8BfJ���|��[����Ω���� F u|g8p��- =����.L��Hy��5����e�.��w"�$`�v�?������6�ss�|A�����#Nfk�Vd�ze�%���?I��d��"���ѓ'O���4������m��u�o�Y�1�����&���w��\h2
���l�����PчQڀ��Ηr� �����D ��%Q�DG��{��d�� ��������y@��	�0���is��*l���� ��s�������� �Ҧ�6_B�����D��0��� �:e����!ϩ<H6`,�Q�싻= l3a+i����6�F���N��2t`���~����[v�(�m<u��������ٕ��1����W����-�hS�G򀍱��>9�
 ����,�h�|� >��U�D@����ɺ�G�g���-G��HK= ���X�7:M�tG����@�&)Y�~���W�^g�^�mp�`�����Jro���L�w�Eg�q�\M��F�3����!`��g���r5����-
��dʉ�\�3a�aa@���BO߾�iV��#kXr�tX�`��&��p����:��K��������=����5o8@��͛������Y���}j,B}�R��SK�ԩI]�hQz:�j����Qa�i�\m�2ԟ��43�C?�����3�@�kj`a��xgz�� @�J���l<	s�-nMd��낟�����b ہ�Z�N?|=&�f0O���t�������j~TQ_�����AJP�(22�a�*���h� �8��SnKg@�t\��x���-)���������"\����ҝ�չ��}�m�?�v Z��ڝ(�422����R��Z��}�Pc�m�����4U��I����^z�Y��[��y�ЫF���?��_z�SY���� 2���x@�#�g�u�~Գ����0%_� l�nD>z	�p��Y���X'꓀�����ߋ�����qgr��8����Sz;[�V1��PDD���([ác�3�Ô��#Nf+1l��r	y<�:)R��yȵD-�8������������~��u}=�'�nC]@��ڮ��3At����:+��Ͷ�����=E^K!	4��@Gձ0�'���>#V���P�=ީ�2X"�(	!,�{>�ٮϣ�s��ʪ?6 ���o򁋡xa�^خ�}g����AxY����%���[֘�z�y�qggg�ݛ�BϦ��4��i�ۏЅ���È���J�8�9���(:=��:�H��ԟwy�t<��y1�h���~&$���,�dBDxLi���繈.�*���:���
M����ƾ� 1@�GZX\�y����~��g'�(a���֜�j�?��7�Z @���������A�T<S�'�fͽ�l˲�k�F�K,qe�X�>y�}c	�>P���pu��e�5�?S��{�X5YD45A��)���۠��R�IzUau��J��|��a�L?[:YD��"} ���?ߚ|
X��N�X�ir*�ô�����>�wg��tx���giŀ|��~���C�3q��o���̸8��������i��	��ęWU��N����\K�H$0�9��ݞ�>d���l���vPЎ,�|$a8�q���SJ�z���������x W68xU;#����P|��$�~rV=��:���=�H
	�K�B���_%�kڰA}7V��u�{�P���-�^�,//Cȧ��:��z�;�z�����ὅ���y�9|�d5�׷G���mb��Z�������Ȭ{w:��s�.�e������
����GbNs=���m�r�e�227ՙ�%�^o�/��Y���4�֦�o�S��(X
�����~7:�!�	v���w�Kr�B��bi��S�$0�����Rw��t��}
1?��9萤��k�,�ֵD���O�X���\��1�q=��mέ�;�#m�Ʒ�j.�\Y!��WWjh�	�?�*�t//'cD"��ͺ���h����#jF�PQܜ�f�������g��ɹ��AY��E���>��D���*.��:�q�Y9�)(萟O�T*�ˬ��X�H�����T|999�Sndd�=�c�8�Tݼ��ې�T��P���»E�7k�ckk�6-�y[X��j�]�l���k���S��%� �XG�oB�P,,�Z�>����rQ���;sE!*��c���[ ��F���8XD������T���[W?�0y����,�T�A��v"�V�A����y�~��ݫi�n�A�N�>��w�l*ܬ��u`��B����j9*��ʢӉ��C� z��;�����D;��=�Fv�`�:��n�O��8�fsN@@ �˽��pdd$�Ϩ����I���''�w�O{��6;��bǖ|n�u_�wq8o�?~FB�]٘��/AdIqqi�����S�}��^��J�Z�ʼ�$�)i�C�L��.���]�_U�02���G��n�0I4^"�|���pSî�4�a��뮏eQߦ�&x$G�]="��M�`"�]��s&����Rͽe�w���G����Xl����w� ���[%��gR�s�dqC7C��������Ph��InI�y2�����-����u{�|b�ǔ4����x��V�:� ��tG����N)�]�&�G�>.
|{NR��Q�5�A�� PK   ��eT����
       jsons/user_defined.json��ۊ�0�_e�u,t�d�4��EKiS(�P|��*^���Ky���&�E��T�53��Hށv[)�]���ʵQX�?�ntil A�]i��Om������1~�k�w�o6'�[�P�[��Z����Y ���\FB
��x�<A�P��P��y�,�s,]�u�N�_�&�u��^d}��L<�̃����7y	�;`�Ǖn�"޾-�?�!���Y/���S�F"$�@�����
�}�����ۮ�	e�{�taWB��]`EQ�Qݼ1�ϲ��Ǎq��|�_�Gc��%t�6q���l����7����>��do��Ru��콖��JG��_����wsL-9�('*�a��0�U�1ayFs)DB=L=U�L����蜫	��C�JWs�`B.0�0��6�>������;�e��>���d��v#_�������Q|�b�}{M���r���x�������ϼ��ޮ�g� qÑ�������vGv����Ў�އ0v���y����}}�7��PK
   ��eT"�e�  ]�                   cirkitFile.jsonPK
   ѕeTד���l  V�  /               images/96360f2e-15f0-4a95-ae8d-a24fd3f977b3.jpgPK
   �beTT�a�f�  ً  /             *|  images/f9879790-346d-4fb7-a00c-c72301b216f4.pngPK
   ��eT����
                 � jsons/user_defined.jsonPK      <  	   